.title Crossbar Circuit
.lib /root/miniforge3/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.subckt mlp NUDGED FREE X_0 X_1 X_2 X_3 Y_0_NUDGED
.subckt synapse WWL WBL RIN ROUT REF
Swrite_nfet MEM WBL WWL 0 switch
Ccap MEM REF 0.05pF capacitor
Xread_nfet RIN MEM ROUT REF sky130_fd_pr__nfet_01v8 l=0.15 w=1.0
.ends synapse

.subckt amp_lin IN OUT
Rshort INN OUT 0.0Ohm
Rmeas IN INN 0.001Ohm
ROUT OUT 0 1000kOhm
.ends amp_lin

.subckt amp_pos IN OUT
Rshort INN OUT 0.0Ohm
Rmeas IN INN 0.001Ohm
ROUT OUT 0 1000kOhm
Vdiol DIOL 0 0.65V
Ddiol DIOL IN diode
.ends amp_pos

.subckt amp_neg IN OUT
Rshort INN OUT 0.0Ohm
Rmeas IN INN 0.001Ohm
ROUT OUT 0 1000kOhm
Vdiou DIOU IN 0.65V
Ddiou DIOU 0 diode
.ends amp_neg

.subckt optimizer WBL FREE NUDGED NUDGED_OUTER UPDATE REF
Bopamp OUT 0 v={max(V(WBL), V(REF)+0.6)*V(NUDGED_OUTER)/1.95}
Sstore OUT STORE NUDGED 0 switch
Cstore STORE 0 0.5pF capacitor
Sread STORE WBL UPDATE 0 switch
.ends optimizer

.subckt crossbar_0 FREE NUDGED NUDGED_OUTER UPDATE RIN_0 RIN_1 RIN_2 RIN_3 ROUT_0 ROUT_1 ROUT_2 ROUT_3 ROUT_4 ROUT_5 ROUT_6 ROUT_7 ROUT_8 ROUT_9 ROUT_10 ROUT_11 ROUT_12 ROUT_13 ROUT_14 ROUT_15
XW_0_0 WWL_0 WBL_0 RIN_0 ROUT_0 REF_0_0 synapse
Rref_0_0 REF_0_0 ROUT_0 0
Sref_0_0 REF_0 REF_0_0 WWL_0 0 switch
XW_0_1 WWL_0 WBL_1 RIN_0 ROUT_1 REF_0_1 synapse
Rref_0_1 REF_0_1 ROUT_1 0
Sref_0_1 REF_1 REF_0_1 WWL_0 0 switch
XW_0_2 WWL_0 WBL_2 RIN_0 ROUT_2 REF_0_2 synapse
Rref_0_2 REF_0_2 ROUT_2 0
Sref_0_2 REF_2 REF_0_2 WWL_0 0 switch
XW_0_3 WWL_0 WBL_3 RIN_0 ROUT_3 REF_0_3 synapse
Rref_0_3 REF_0_3 ROUT_3 0
Sref_0_3 REF_3 REF_0_3 WWL_0 0 switch
XW_0_4 WWL_0 WBL_4 RIN_0 ROUT_4 REF_0_4 synapse
Rref_0_4 REF_0_4 ROUT_4 0
Sref_0_4 REF_4 REF_0_4 WWL_0 0 switch
XW_0_5 WWL_0 WBL_5 RIN_0 ROUT_5 REF_0_5 synapse
Rref_0_5 REF_0_5 ROUT_5 0
Sref_0_5 REF_5 REF_0_5 WWL_0 0 switch
XW_0_6 WWL_0 WBL_6 RIN_0 ROUT_6 REF_0_6 synapse
Rref_0_6 REF_0_6 ROUT_6 0
Sref_0_6 REF_6 REF_0_6 WWL_0 0 switch
XW_0_7 WWL_0 WBL_7 RIN_0 ROUT_7 REF_0_7 synapse
Rref_0_7 REF_0_7 ROUT_7 0
Sref_0_7 REF_7 REF_0_7 WWL_0 0 switch
XW_0_8 WWL_0 WBL_8 RIN_0 ROUT_8 REF_0_8 synapse
Rref_0_8 REF_0_8 ROUT_8 0
Sref_0_8 REF_8 REF_0_8 WWL_0 0 switch
XW_0_9 WWL_0 WBL_9 RIN_0 ROUT_9 REF_0_9 synapse
Rref_0_9 REF_0_9 ROUT_9 0
Sref_0_9 REF_9 REF_0_9 WWL_0 0 switch
XW_0_10 WWL_0 WBL_10 RIN_0 ROUT_10 REF_0_10 synapse
Rref_0_10 REF_0_10 ROUT_10 0
Sref_0_10 REF_10 REF_0_10 WWL_0 0 switch
XW_0_11 WWL_0 WBL_11 RIN_0 ROUT_11 REF_0_11 synapse
Rref_0_11 REF_0_11 ROUT_11 0
Sref_0_11 REF_11 REF_0_11 WWL_0 0 switch
XW_0_12 WWL_0 WBL_12 RIN_0 ROUT_12 REF_0_12 synapse
Rref_0_12 REF_0_12 ROUT_12 0
Sref_0_12 REF_12 REF_0_12 WWL_0 0 switch
XW_0_13 WWL_0 WBL_13 RIN_0 ROUT_13 REF_0_13 synapse
Rref_0_13 REF_0_13 ROUT_13 0
Sref_0_13 REF_13 REF_0_13 WWL_0 0 switch
XW_0_14 WWL_0 WBL_14 RIN_0 ROUT_14 REF_0_14 synapse
Rref_0_14 REF_0_14 ROUT_14 0
Sref_0_14 REF_14 REF_0_14 WWL_0 0 switch
XW_0_15 WWL_0 WBL_15 RIN_0 ROUT_15 REF_0_15 synapse
Rref_0_15 REF_0_15 ROUT_15 0
Sref_0_15 REF_15 REF_0_15 WWL_0 0 switch
XW_1_0 WWL_1 WBL_0 RIN_1 ROUT_0 REF_1_0 synapse
Rref_1_0 REF_1_0 ROUT_0 0
Sref_1_0 REF_0 REF_1_0 WWL_1 0 switch
XW_1_1 WWL_1 WBL_1 RIN_1 ROUT_1 REF_1_1 synapse
Rref_1_1 REF_1_1 ROUT_1 0
Sref_1_1 REF_1 REF_1_1 WWL_1 0 switch
XW_1_2 WWL_1 WBL_2 RIN_1 ROUT_2 REF_1_2 synapse
Rref_1_2 REF_1_2 ROUT_2 0
Sref_1_2 REF_2 REF_1_2 WWL_1 0 switch
XW_1_3 WWL_1 WBL_3 RIN_1 ROUT_3 REF_1_3 synapse
Rref_1_3 REF_1_3 ROUT_3 0
Sref_1_3 REF_3 REF_1_3 WWL_1 0 switch
XW_1_4 WWL_1 WBL_4 RIN_1 ROUT_4 REF_1_4 synapse
Rref_1_4 REF_1_4 ROUT_4 0
Sref_1_4 REF_4 REF_1_4 WWL_1 0 switch
XW_1_5 WWL_1 WBL_5 RIN_1 ROUT_5 REF_1_5 synapse
Rref_1_5 REF_1_5 ROUT_5 0
Sref_1_5 REF_5 REF_1_5 WWL_1 0 switch
XW_1_6 WWL_1 WBL_6 RIN_1 ROUT_6 REF_1_6 synapse
Rref_1_6 REF_1_6 ROUT_6 0
Sref_1_6 REF_6 REF_1_6 WWL_1 0 switch
XW_1_7 WWL_1 WBL_7 RIN_1 ROUT_7 REF_1_7 synapse
Rref_1_7 REF_1_7 ROUT_7 0
Sref_1_7 REF_7 REF_1_7 WWL_1 0 switch
XW_1_8 WWL_1 WBL_8 RIN_1 ROUT_8 REF_1_8 synapse
Rref_1_8 REF_1_8 ROUT_8 0
Sref_1_8 REF_8 REF_1_8 WWL_1 0 switch
XW_1_9 WWL_1 WBL_9 RIN_1 ROUT_9 REF_1_9 synapse
Rref_1_9 REF_1_9 ROUT_9 0
Sref_1_9 REF_9 REF_1_9 WWL_1 0 switch
XW_1_10 WWL_1 WBL_10 RIN_1 ROUT_10 REF_1_10 synapse
Rref_1_10 REF_1_10 ROUT_10 0
Sref_1_10 REF_10 REF_1_10 WWL_1 0 switch
XW_1_11 WWL_1 WBL_11 RIN_1 ROUT_11 REF_1_11 synapse
Rref_1_11 REF_1_11 ROUT_11 0
Sref_1_11 REF_11 REF_1_11 WWL_1 0 switch
XW_1_12 WWL_1 WBL_12 RIN_1 ROUT_12 REF_1_12 synapse
Rref_1_12 REF_1_12 ROUT_12 0
Sref_1_12 REF_12 REF_1_12 WWL_1 0 switch
XW_1_13 WWL_1 WBL_13 RIN_1 ROUT_13 REF_1_13 synapse
Rref_1_13 REF_1_13 ROUT_13 0
Sref_1_13 REF_13 REF_1_13 WWL_1 0 switch
XW_1_14 WWL_1 WBL_14 RIN_1 ROUT_14 REF_1_14 synapse
Rref_1_14 REF_1_14 ROUT_14 0
Sref_1_14 REF_14 REF_1_14 WWL_1 0 switch
XW_1_15 WWL_1 WBL_15 RIN_1 ROUT_15 REF_1_15 synapse
Rref_1_15 REF_1_15 ROUT_15 0
Sref_1_15 REF_15 REF_1_15 WWL_1 0 switch
XW_2_0 WWL_2 WBL_0 RIN_2 ROUT_0 REF_2_0 synapse
Rref_2_0 REF_2_0 ROUT_0 0
Sref_2_0 REF_0 REF_2_0 WWL_2 0 switch
XW_2_1 WWL_2 WBL_1 RIN_2 ROUT_1 REF_2_1 synapse
Rref_2_1 REF_2_1 ROUT_1 0
Sref_2_1 REF_1 REF_2_1 WWL_2 0 switch
XW_2_2 WWL_2 WBL_2 RIN_2 ROUT_2 REF_2_2 synapse
Rref_2_2 REF_2_2 ROUT_2 0
Sref_2_2 REF_2 REF_2_2 WWL_2 0 switch
XW_2_3 WWL_2 WBL_3 RIN_2 ROUT_3 REF_2_3 synapse
Rref_2_3 REF_2_3 ROUT_3 0
Sref_2_3 REF_3 REF_2_3 WWL_2 0 switch
XW_2_4 WWL_2 WBL_4 RIN_2 ROUT_4 REF_2_4 synapse
Rref_2_4 REF_2_4 ROUT_4 0
Sref_2_4 REF_4 REF_2_4 WWL_2 0 switch
XW_2_5 WWL_2 WBL_5 RIN_2 ROUT_5 REF_2_5 synapse
Rref_2_5 REF_2_5 ROUT_5 0
Sref_2_5 REF_5 REF_2_5 WWL_2 0 switch
XW_2_6 WWL_2 WBL_6 RIN_2 ROUT_6 REF_2_6 synapse
Rref_2_6 REF_2_6 ROUT_6 0
Sref_2_6 REF_6 REF_2_6 WWL_2 0 switch
XW_2_7 WWL_2 WBL_7 RIN_2 ROUT_7 REF_2_7 synapse
Rref_2_7 REF_2_7 ROUT_7 0
Sref_2_7 REF_7 REF_2_7 WWL_2 0 switch
XW_2_8 WWL_2 WBL_8 RIN_2 ROUT_8 REF_2_8 synapse
Rref_2_8 REF_2_8 ROUT_8 0
Sref_2_8 REF_8 REF_2_8 WWL_2 0 switch
XW_2_9 WWL_2 WBL_9 RIN_2 ROUT_9 REF_2_9 synapse
Rref_2_9 REF_2_9 ROUT_9 0
Sref_2_9 REF_9 REF_2_9 WWL_2 0 switch
XW_2_10 WWL_2 WBL_10 RIN_2 ROUT_10 REF_2_10 synapse
Rref_2_10 REF_2_10 ROUT_10 0
Sref_2_10 REF_10 REF_2_10 WWL_2 0 switch
XW_2_11 WWL_2 WBL_11 RIN_2 ROUT_11 REF_2_11 synapse
Rref_2_11 REF_2_11 ROUT_11 0
Sref_2_11 REF_11 REF_2_11 WWL_2 0 switch
XW_2_12 WWL_2 WBL_12 RIN_2 ROUT_12 REF_2_12 synapse
Rref_2_12 REF_2_12 ROUT_12 0
Sref_2_12 REF_12 REF_2_12 WWL_2 0 switch
XW_2_13 WWL_2 WBL_13 RIN_2 ROUT_13 REF_2_13 synapse
Rref_2_13 REF_2_13 ROUT_13 0
Sref_2_13 REF_13 REF_2_13 WWL_2 0 switch
XW_2_14 WWL_2 WBL_14 RIN_2 ROUT_14 REF_2_14 synapse
Rref_2_14 REF_2_14 ROUT_14 0
Sref_2_14 REF_14 REF_2_14 WWL_2 0 switch
XW_2_15 WWL_2 WBL_15 RIN_2 ROUT_15 REF_2_15 synapse
Rref_2_15 REF_2_15 ROUT_15 0
Sref_2_15 REF_15 REF_2_15 WWL_2 0 switch
XW_3_0 WWL_3 WBL_0 RIN_3 ROUT_0 REF_3_0 synapse
Rref_3_0 REF_3_0 ROUT_0 0
Sref_3_0 REF_0 REF_3_0 WWL_3 0 switch
XW_3_1 WWL_3 WBL_1 RIN_3 ROUT_1 REF_3_1 synapse
Rref_3_1 REF_3_1 ROUT_1 0
Sref_3_1 REF_1 REF_3_1 WWL_3 0 switch
XW_3_2 WWL_3 WBL_2 RIN_3 ROUT_2 REF_3_2 synapse
Rref_3_2 REF_3_2 ROUT_2 0
Sref_3_2 REF_2 REF_3_2 WWL_3 0 switch
XW_3_3 WWL_3 WBL_3 RIN_3 ROUT_3 REF_3_3 synapse
Rref_3_3 REF_3_3 ROUT_3 0
Sref_3_3 REF_3 REF_3_3 WWL_3 0 switch
XW_3_4 WWL_3 WBL_4 RIN_3 ROUT_4 REF_3_4 synapse
Rref_3_4 REF_3_4 ROUT_4 0
Sref_3_4 REF_4 REF_3_4 WWL_3 0 switch
XW_3_5 WWL_3 WBL_5 RIN_3 ROUT_5 REF_3_5 synapse
Rref_3_5 REF_3_5 ROUT_5 0
Sref_3_5 REF_5 REF_3_5 WWL_3 0 switch
XW_3_6 WWL_3 WBL_6 RIN_3 ROUT_6 REF_3_6 synapse
Rref_3_6 REF_3_6 ROUT_6 0
Sref_3_6 REF_6 REF_3_6 WWL_3 0 switch
XW_3_7 WWL_3 WBL_7 RIN_3 ROUT_7 REF_3_7 synapse
Rref_3_7 REF_3_7 ROUT_7 0
Sref_3_7 REF_7 REF_3_7 WWL_3 0 switch
XW_3_8 WWL_3 WBL_8 RIN_3 ROUT_8 REF_3_8 synapse
Rref_3_8 REF_3_8 ROUT_8 0
Sref_3_8 REF_8 REF_3_8 WWL_3 0 switch
XW_3_9 WWL_3 WBL_9 RIN_3 ROUT_9 REF_3_9 synapse
Rref_3_9 REF_3_9 ROUT_9 0
Sref_3_9 REF_9 REF_3_9 WWL_3 0 switch
XW_3_10 WWL_3 WBL_10 RIN_3 ROUT_10 REF_3_10 synapse
Rref_3_10 REF_3_10 ROUT_10 0
Sref_3_10 REF_10 REF_3_10 WWL_3 0 switch
XW_3_11 WWL_3 WBL_11 RIN_3 ROUT_11 REF_3_11 synapse
Rref_3_11 REF_3_11 ROUT_11 0
Sref_3_11 REF_11 REF_3_11 WWL_3 0 switch
XW_3_12 WWL_3 WBL_12 RIN_3 ROUT_12 REF_3_12 synapse
Rref_3_12 REF_3_12 ROUT_12 0
Sref_3_12 REF_12 REF_3_12 WWL_3 0 switch
XW_3_13 WWL_3 WBL_13 RIN_3 ROUT_13 REF_3_13 synapse
Rref_3_13 REF_3_13 ROUT_13 0
Sref_3_13 REF_13 REF_3_13 WWL_3 0 switch
XW_3_14 WWL_3 WBL_14 RIN_3 ROUT_14 REF_3_14 synapse
Rref_3_14 REF_3_14 ROUT_14 0
Sref_3_14 REF_14 REF_3_14 WWL_3 0 switch
XW_3_15 WWL_3 WBL_15 RIN_3 ROUT_15 REF_3_15 synapse
Rref_3_15 REF_3_15 ROUT_15 0
Sref_3_15 REF_15 REF_3_15 WWL_3 0 switch
Xopt_0 WBL_0 FREE NUDGED NUDGED_OUTER UPDATE REF_0 optimizer
SGND_0 REF_0 0 SET 0 switch
Xopt_1 WBL_1 FREE NUDGED NUDGED_OUTER UPDATE REF_1 optimizer
SGND_1 REF_1 0 SET 0 switch
Xopt_2 WBL_2 FREE NUDGED NUDGED_OUTER UPDATE REF_2 optimizer
SGND_2 REF_2 0 SET 0 switch
Xopt_3 WBL_3 FREE NUDGED NUDGED_OUTER UPDATE REF_3 optimizer
SGND_3 REF_3 0 SET 0 switch
Xopt_4 WBL_4 FREE NUDGED NUDGED_OUTER UPDATE REF_4 optimizer
SGND_4 REF_4 0 SET 0 switch
Xopt_5 WBL_5 FREE NUDGED NUDGED_OUTER UPDATE REF_5 optimizer
SGND_5 REF_5 0 SET 0 switch
Xopt_6 WBL_6 FREE NUDGED NUDGED_OUTER UPDATE REF_6 optimizer
SGND_6 REF_6 0 SET 0 switch
Xopt_7 WBL_7 FREE NUDGED NUDGED_OUTER UPDATE REF_7 optimizer
SGND_7 REF_7 0 SET 0 switch
Xopt_8 WBL_8 FREE NUDGED NUDGED_OUTER UPDATE REF_8 optimizer
SGND_8 REF_8 0 SET 0 switch
Xopt_9 WBL_9 FREE NUDGED NUDGED_OUTER UPDATE REF_9 optimizer
SGND_9 REF_9 0 SET 0 switch
Xopt_10 WBL_10 FREE NUDGED NUDGED_OUTER UPDATE REF_10 optimizer
SGND_10 REF_10 0 SET 0 switch
Xopt_11 WBL_11 FREE NUDGED NUDGED_OUTER UPDATE REF_11 optimizer
SGND_11 REF_11 0 SET 0 switch
Xopt_12 WBL_12 FREE NUDGED NUDGED_OUTER UPDATE REF_12 optimizer
SGND_12 REF_12 0 SET 0 switch
Xopt_13 WBL_13 FREE NUDGED NUDGED_OUTER UPDATE REF_13 optimizer
SGND_13 REF_13 0 SET 0 switch
Xopt_14 WBL_14 FREE NUDGED NUDGED_OUTER UPDATE REF_14 optimizer
SGND_14 REF_14 0 SET 0 switch
Xopt_15 WBL_15 FREE NUDGED NUDGED_OUTER UPDATE REF_15 optimizer
SGND_15 REF_15 0 SET 0 switch
VSET_0 SET_0 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 0.9829480051994324V 2560.0ns 0.9829480051994324V 2600.0ns 0V 3040.0ns 0V 3080.0ns 2.080735683441162V 4160.0ns 2.080735683441162V 4200.0ns 0V 4640.0ns 0V 4680.0ns 0.9873619675636292V 5760.0ns 0.9873619675636292V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.0302115678787231V 7360.0ns 1.0302115678787231V 7400.0ns 0V)
SSET_0 SET_0 WBL_0 SET 0 switch
VSET_1 SET_1 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.2108234167099V 2560.0ns 1.2108234167099V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.3977434635162354V 4160.0ns 1.3977434635162354V 4200.0ns 0V 4640.0ns 0V 4680.0ns 0.7828106880187988V 5760.0ns 0.7828106880187988V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.0384502410888672V 7360.0ns 1.0384502410888672V 7400.0ns 0V)
SSET_1 SET_1 WBL_1 SET 0 switch
VSET_2 SET_2 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.8060978651046753V 2560.0ns 1.8060978651046753V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.3326979875564575V 4160.0ns 1.3326979875564575V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.910875916481018V 5760.0ns 1.910875916481018V 5800.0ns 0V 6240.0ns 0V 6280.0ns 0.8942763209342957V 7360.0ns 0.8942763209342957V 7400.0ns 0V)
SSET_2 SET_2 WBL_2 SET 0 switch
VSET_3 SET_3 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.329432725906372V 2560.0ns 1.329432725906372V 2600.0ns 0V 3040.0ns 0V 3080.0ns 0.6986654996871948V 4160.0ns 0.6986654996871948V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.0864973068237305V 5760.0ns 1.0864973068237305V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.9976892471313477V 7360.0ns 1.9976892471313477V 7400.0ns 0V)
SSET_3 SET_3 WBL_3 SET 0 switch
VSET_4 SET_4 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 0.8341853022575378V 2560.0ns 0.8341853022575378V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.9504483938217163V 4160.0ns 1.9504483938217163V 4200.0ns 0V 4640.0ns 0V 4680.0ns 0.8567845225334167V 5760.0ns 0.8567845225334167V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.582169771194458V 7360.0ns 1.582169771194458V 7400.0ns 0V)
SSET_4 SET_4 WBL_4 SET 0 switch
VSET_5 SET_5 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.5533759593963623V 2560.0ns 1.5533759593963623V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.81326162815094V 4160.0ns 1.81326162815094V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.332613468170166V 5760.0ns 1.332613468170166V 5800.0ns 0V 6240.0ns 0V 6280.0ns 2.062844753265381V 7360.0ns 2.062844753265381V 7400.0ns 0V)
SSET_5 SET_5 WBL_5 SET 0 switch
VSET_6 SET_6 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.8792916536331177V 2560.0ns 1.8792916536331177V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.0399619340896606V 4160.0ns 1.0399619340896606V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.7082468271255493V 5760.0ns 1.7082468271255493V 5800.0ns 0V 6240.0ns 0V 6280.0ns 2.133021593093872V 7360.0ns 2.133021593093872V 7400.0ns 0V)
SSET_6 SET_6 WBL_6 SET 0 switch
VSET_7 SET_7 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.6415224075317383V 2560.0ns 1.6415224075317383V 2600.0ns 0V 3040.0ns 0V 3080.0ns 0.6575799584388733V 4160.0ns 0.6575799584388733V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.5319570302963257V 5760.0ns 1.5319570302963257V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.6667371988296509V 7360.0ns 1.6667371988296509V 7400.0ns 0V)
SSET_7 SET_7 WBL_7 SET 0 switch
VSET_8 SET_8 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.5379269123077393V 2560.0ns 1.5379269123077393V 2600.0ns 0V 3040.0ns 0V 3080.0ns 0.8200723528862V 4160.0ns 0.8200723528862V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.4644289016723633V 5760.0ns 1.4644289016723633V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.4344080686569214V 7360.0ns 1.4344080686569214V 7400.0ns 0V)
SSET_8 SET_8 WBL_8 SET 0 switch
VSET_9 SET_9 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 2.25247859954834V 2560.0ns 2.25247859954834V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.0413131713867188V 4160.0ns 1.0413131713867188V 4200.0ns 0V 4640.0ns 0V 4680.0ns 2.2179665565490723V 5760.0ns 2.2179665565490723V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.0393548011779785V 7360.0ns 1.0393548011779785V 7400.0ns 0V)
SSET_9 SET_9 WBL_9 SET 0 switch
VSET_10 SET_10 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.4690637588500977V 2560.0ns 1.4690637588500977V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.8613654375076294V 4160.0ns 1.8613654375076294V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.205824613571167V 5760.0ns 1.205824613571167V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.1166459321975708V 7360.0ns 1.1166459321975708V 7400.0ns 0V)
SSET_10 SET_10 WBL_10 SET 0 switch
VSET_11 SET_11 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.281296968460083V 2560.0ns 1.281296968460083V 2600.0ns 0V 3040.0ns 0V 3080.0ns 0.6113315224647522V 4160.0ns 0.6113315224647522V 4200.0ns 0V 4640.0ns 0V 4680.0ns 1.494778037071228V 5760.0ns 1.494778037071228V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.7445769309997559V 7360.0ns 1.7445769309997559V 7400.0ns 0V)
SSET_11 SET_11 WBL_11 SET 0 switch
VSET_12 SET_12 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 2.3497495651245117V 2560.0ns 2.3497495651245117V 2600.0ns 0V 3040.0ns 0V 3080.0ns 0.8706896305084229V 4160.0ns 0.8706896305084229V 4200.0ns 0V 4640.0ns 0V 4680.0ns 2.2397103309631348V 5760.0ns 2.2397103309631348V 5800.0ns 0V 6240.0ns 0V 6280.0ns 2.0292301177978516V 7360.0ns 2.0292301177978516V 7400.0ns 0V)
SSET_12 SET_12 WBL_12 SET 0 switch
VSET_13 SET_13 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 0.7101213335990906V 2560.0ns 0.7101213335990906V 2600.0ns 0V 3040.0ns 0V 3080.0ns 2.1259000301361084V 4160.0ns 2.1259000301361084V 4200.0ns 0V 4640.0ns 0V 4680.0ns 0.8567798137664795V 5760.0ns 0.8567798137664795V 5800.0ns 0V 6240.0ns 0V 6280.0ns 2.3535304069519043V 7360.0ns 2.3535304069519043V 7400.0ns 0V)
SSET_13 SET_13 WBL_13 SET 0 switch
VSET_14 SET_14 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.3132052421569824V 2560.0ns 1.3132052421569824V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.5909745693206787V 4160.0ns 1.5909745693206787V 4200.0ns 0V 4640.0ns 0V 4680.0ns 0.9934470653533936V 5760.0ns 0.9934470653533936V 5800.0ns 0V 6240.0ns 0V 6280.0ns 1.1073631048202515V 7360.0ns 1.1073631048202515V 7400.0ns 0V)
SSET_14 SET_14 WBL_14 SET 0 switch
VSET_15 SET_15 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.501501202583313V 2560.0ns 1.501501202583313V 2600.0ns 0V 3040.0ns 0V 3080.0ns 1.9817596673965454V 4160.0ns 1.9817596673965454V 4200.0ns 0V 4640.0ns 0V 4680.0ns 2.1967568397521973V 5760.0ns 2.1967568397521973V 5800.0ns 0V 6240.0ns 0V 6280.0ns 0.9888023138046265V 7360.0ns 0.9888023138046265V 7400.0ns 0V)
SSET_15 SET_15 WBL_15 SET 0 switch
VSET SET 0 PWL(0ns 1.95V 8000.0ns 1.95V 8040.0ns 0V)
VWWL_0 WWL_0 0 PWL(0ns 0V 1600.0ns 0V 1640.0ns 1.95V 2400.0ns 1.95V 2440.0ns 0V 9600.0ns 0V)
VWWL_1 WWL_1 0 PWL(0ns 0V 3200.0ns 0V 3240.0ns 1.95V 4000.0ns 1.95V 4040.0ns 0V 9600.0ns 0V)
VWWL_2 WWL_2 0 PWL(0ns 0V 4800.0ns 0V 4840.0ns 1.95V 5600.0ns 1.95V 5640.0ns 0V 9600.0ns 0V)
VWWL_3 WWL_3 0 PWL(0ns 0V 6400.0ns 0V 6440.0ns 1.95V 7200.0ns 1.95V 7240.0ns 0V 9600.0ns 0V)
.ends crossbar_0

.subckt crossbar_1 FREE NUDGED NUDGED_OUTER UPDATE RIN_0 RIN_1 RIN_2 RIN_3 RIN_4 RIN_5 RIN_6 RIN_7 RIN_8 RIN_9 RIN_10 RIN_11 RIN_12 RIN_13 RIN_14 RIN_15 ROUT_0
XW_0_0 WWL_0 WBL_0 RIN_0 ROUT_0 REF_0_0 synapse
Rref_0_0 REF_0_0 ROUT_0 0
Sref_0_0 REF_0 REF_0_0 WWL_0 0 switch
XW_1_0 WWL_0 WBL_1 RIN_1 ROUT_0 REF_1_0 synapse
Rref_1_0 REF_1_0 ROUT_0 0
Sref_1_0 REF_1 REF_1_0 WWL_0 0 switch
XW_2_0 WWL_0 WBL_2 RIN_2 ROUT_0 REF_2_0 synapse
Rref_2_0 REF_2_0 ROUT_0 0
Sref_2_0 REF_2 REF_2_0 WWL_0 0 switch
XW_3_0 WWL_0 WBL_3 RIN_3 ROUT_0 REF_3_0 synapse
Rref_3_0 REF_3_0 ROUT_0 0
Sref_3_0 REF_3 REF_3_0 WWL_0 0 switch
XW_4_0 WWL_0 WBL_4 RIN_4 ROUT_0 REF_4_0 synapse
Rref_4_0 REF_4_0 ROUT_0 0
Sref_4_0 REF_4 REF_4_0 WWL_0 0 switch
XW_5_0 WWL_0 WBL_5 RIN_5 ROUT_0 REF_5_0 synapse
Rref_5_0 REF_5_0 ROUT_0 0
Sref_5_0 REF_5 REF_5_0 WWL_0 0 switch
XW_6_0 WWL_0 WBL_6 RIN_6 ROUT_0 REF_6_0 synapse
Rref_6_0 REF_6_0 ROUT_0 0
Sref_6_0 REF_6 REF_6_0 WWL_0 0 switch
XW_7_0 WWL_0 WBL_7 RIN_7 ROUT_0 REF_7_0 synapse
Rref_7_0 REF_7_0 ROUT_0 0
Sref_7_0 REF_7 REF_7_0 WWL_0 0 switch
XW_8_0 WWL_0 WBL_8 RIN_8 ROUT_0 REF_8_0 synapse
Rref_8_0 REF_8_0 ROUT_0 0
Sref_8_0 REF_8 REF_8_0 WWL_0 0 switch
XW_9_0 WWL_0 WBL_9 RIN_9 ROUT_0 REF_9_0 synapse
Rref_9_0 REF_9_0 ROUT_0 0
Sref_9_0 REF_9 REF_9_0 WWL_0 0 switch
XW_10_0 WWL_0 WBL_10 RIN_10 ROUT_0 REF_10_0 synapse
Rref_10_0 REF_10_0 ROUT_0 0
Sref_10_0 REF_10 REF_10_0 WWL_0 0 switch
XW_11_0 WWL_0 WBL_11 RIN_11 ROUT_0 REF_11_0 synapse
Rref_11_0 REF_11_0 ROUT_0 0
Sref_11_0 REF_11 REF_11_0 WWL_0 0 switch
XW_12_0 WWL_0 WBL_12 RIN_12 ROUT_0 REF_12_0 synapse
Rref_12_0 REF_12_0 ROUT_0 0
Sref_12_0 REF_12 REF_12_0 WWL_0 0 switch
XW_13_0 WWL_0 WBL_13 RIN_13 ROUT_0 REF_13_0 synapse
Rref_13_0 REF_13_0 ROUT_0 0
Sref_13_0 REF_13 REF_13_0 WWL_0 0 switch
XW_14_0 WWL_0 WBL_14 RIN_14 ROUT_0 REF_14_0 synapse
Rref_14_0 REF_14_0 ROUT_0 0
Sref_14_0 REF_14 REF_14_0 WWL_0 0 switch
XW_15_0 WWL_0 WBL_15 RIN_15 ROUT_0 REF_15_0 synapse
Rref_15_0 REF_15_0 ROUT_0 0
Sref_15_0 REF_15 REF_15_0 WWL_0 0 switch
Xopt_0 WBL_0 FREE NUDGED NUDGED_OUTER UPDATE REF_0 optimizer
SGND_0 REF_0 0 SET 0 switch
Xopt_1 WBL_1 FREE NUDGED NUDGED_OUTER UPDATE REF_1 optimizer
SGND_1 REF_1 0 SET 0 switch
Xopt_2 WBL_2 FREE NUDGED NUDGED_OUTER UPDATE REF_2 optimizer
SGND_2 REF_2 0 SET 0 switch
Xopt_3 WBL_3 FREE NUDGED NUDGED_OUTER UPDATE REF_3 optimizer
SGND_3 REF_3 0 SET 0 switch
Xopt_4 WBL_4 FREE NUDGED NUDGED_OUTER UPDATE REF_4 optimizer
SGND_4 REF_4 0 SET 0 switch
Xopt_5 WBL_5 FREE NUDGED NUDGED_OUTER UPDATE REF_5 optimizer
SGND_5 REF_5 0 SET 0 switch
Xopt_6 WBL_6 FREE NUDGED NUDGED_OUTER UPDATE REF_6 optimizer
SGND_6 REF_6 0 SET 0 switch
Xopt_7 WBL_7 FREE NUDGED NUDGED_OUTER UPDATE REF_7 optimizer
SGND_7 REF_7 0 SET 0 switch
Xopt_8 WBL_8 FREE NUDGED NUDGED_OUTER UPDATE REF_8 optimizer
SGND_8 REF_8 0 SET 0 switch
Xopt_9 WBL_9 FREE NUDGED NUDGED_OUTER UPDATE REF_9 optimizer
SGND_9 REF_9 0 SET 0 switch
Xopt_10 WBL_10 FREE NUDGED NUDGED_OUTER UPDATE REF_10 optimizer
SGND_10 REF_10 0 SET 0 switch
Xopt_11 WBL_11 FREE NUDGED NUDGED_OUTER UPDATE REF_11 optimizer
SGND_11 REF_11 0 SET 0 switch
Xopt_12 WBL_12 FREE NUDGED NUDGED_OUTER UPDATE REF_12 optimizer
SGND_12 REF_12 0 SET 0 switch
Xopt_13 WBL_13 FREE NUDGED NUDGED_OUTER UPDATE REF_13 optimizer
SGND_13 REF_13 0 SET 0 switch
Xopt_14 WBL_14 FREE NUDGED NUDGED_OUTER UPDATE REF_14 optimizer
SGND_14 REF_14 0 SET 0 switch
Xopt_15 WBL_15 FREE NUDGED NUDGED_OUTER UPDATE REF_15 optimizer
SGND_15 REF_15 0 SET 0 switch
VSET_0 SET_0 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 2.2431302070617676V 2560.0ns 2.2431302070617676V 2600.0ns 0V)
SSET_0 SET_0 WBL_0 SET 0 switch
VSET_1 SET_1 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 0.8953609466552734V 2560.0ns 0.8953609466552734V 2600.0ns 0V)
SSET_1 SET_1 WBL_1 SET 0 switch
VSET_2 SET_2 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.9847131967544556V 2560.0ns 1.9847131967544556V 2600.0ns 0V)
SSET_2 SET_2 WBL_2 SET 0 switch
VSET_3 SET_3 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.1838825941085815V 2560.0ns 1.1838825941085815V 2600.0ns 0V)
SSET_3 SET_3 WBL_3 SET 0 switch
VSET_4 SET_4 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 0.6845744848251343V 2560.0ns 0.6845744848251343V 2600.0ns 0V)
SSET_4 SET_4 WBL_4 SET 0 switch
VSET_5 SET_5 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 2.378915786743164V 2560.0ns 2.378915786743164V 2600.0ns 0V)
SSET_5 SET_5 WBL_5 SET 0 switch
VSET_6 SET_6 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 0.6850359439849854V 2560.0ns 0.6850359439849854V 2600.0ns 0V)
SSET_6 SET_6 WBL_6 SET 0 switch
VSET_7 SET_7 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 2.2427480220794678V 2560.0ns 2.2427480220794678V 2600.0ns 0V)
SSET_7 SET_7 WBL_7 SET 0 switch
VSET_8 SET_8 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 2.011002540588379V 2560.0ns 2.011002540588379V 2600.0ns 0V)
SSET_8 SET_8 WBL_8 SET 0 switch
VSET_9 SET_9 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 2.109861135482788V 2560.0ns 2.109861135482788V 2600.0ns 0V)
SSET_9 SET_9 WBL_9 SET 0 switch
VSET_10 SET_10 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.8774642944335938V 2560.0ns 1.8774642944335938V 2600.0ns 0V)
SSET_10 SET_10 WBL_10 SET 0 switch
VSET_11 SET_11 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.8260143995285034V 2560.0ns 1.8260143995285034V 2600.0ns 0V)
SSET_11 SET_11 WBL_11 SET 0 switch
VSET_12 SET_12 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.6543604135513306V 2560.0ns 1.6543604135513306V 2600.0ns 0V)
SSET_12 SET_12 WBL_12 SET 0 switch
VSET_13 SET_13 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 0.7271312475204468V 2560.0ns 0.7271312475204468V 2600.0ns 0V)
SSET_13 SET_13 WBL_13 SET 0 switch
VSET_14 SET_14 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.3233263492584229V 2560.0ns 1.3233263492584229V 2600.0ns 0V)
SSET_14 SET_14 WBL_14 SET 0 switch
VSET_15 SET_15 0 PWL(0ns 0V 1440.0ns 0V 1480.0ns 1.6358261108398438V 2560.0ns 1.6358261108398438V 2600.0ns 0V)
SSET_15 SET_15 WBL_15 SET 0 switch
VSET SET 0 PWL(0ns 1.95V 8000.0ns 1.95V 8040.0ns 0V)
VWWL_0 WWL_0 0 PWL(0ns 0V 1600.0ns 0V 1640.0ns 1.95V 2400.0ns 1.95V 2440.0ns 0V 9600.0ns 0V)
.ends crossbar_1

.subckt loss FREE NUDGED Y_0 PRED_0
SPRED_0_NUDGED PRED_0 PRED_0_NUDGED NUDGED 0 switch
SPRED_0_FREE PRED_0 PRED_0_FREE FREE 0 switch
CPRED_0_FREE PRED_0_FREE 0 0.05pF capacitor
BNUDGE_0 PRED_0_NUDGED 0 i={-0.001 * (V(Y_0)-V(PRED_0_FREE)) * V(NUDGED)}
BLOSS LOSS 0 v={(V(Y_0)-V(PRED_0))*(V(Y_0)-V(PRED_0))}
.ends loss
Xact_1_0 preact_1_0 postact_1_0 amp_pos
Xact_1_1 preact_1_1 postact_1_1 amp_pos
Xact_1_2 preact_1_2 postact_1_2 amp_pos
Xact_1_3 preact_1_3 postact_1_3 amp_pos
Xact_1_4 preact_1_4 postact_1_4 amp_pos
Xact_1_5 preact_1_5 postact_1_5 amp_pos
Xact_1_6 preact_1_6 postact_1_6 amp_pos
Xact_1_7 preact_1_7 postact_1_7 amp_pos
Xact_1_8 preact_1_8 postact_1_8 amp_pos
Xact_1_9 preact_1_9 postact_1_9 amp_pos
Xact_1_10 preact_1_10 postact_1_10 amp_pos
Xact_1_11 preact_1_11 postact_1_11 amp_pos
Xact_1_12 preact_1_12 postact_1_12 amp_pos
Xact_1_13 preact_1_13 postact_1_13 amp_pos
Xact_1_14 preact_1_14 postact_1_14 amp_pos
Xact_1_15 preact_1_15 postact_1_15 amp_pos
Xact_2_0 preact_2_0 postact_2_0 amp_lin
Xloss FREE NUDGED_OUTER Y_0 postact_2_0 loss
VFREE FREE 0 PWL(0ns 0V 9600.0ns 0V)
VNUDGED NUDGED 0 PWL(0ns 0V 9600.0ns 0V)
VNUDGED_OUTER NUDGED_OUTER 0 PWL(0ns 0V 9600.0ns 0V)
VUPDATE UPDATE 0 PWL(0ns 0V 9600.0ns 0V)
VX_0 postact_0_0 0 PWL(0ns 0V 9600.0ns 0V)
VXn_0 0 postact_0_1 PWL(0ns 0V 9600.0ns 0V)
VX_1 postact_0_2 0 PWL(0ns 0V 9600.0ns 0V)
VXn_1 0 postact_0_3 PWL(0ns 0V 9600.0ns 0V)
VY_0 Y_0 0 PWL(0ns 0V 9600.0ns 0V)
.model switch VSWITCH (ROFF=100000000000.0kOhm RON=0.0001Ohm VOFF=0.4V VON=0.5V)
.model diode D ()
.model capacitor C ()
.ends mlp
Xmlp NUDGED FREE X_0 X_1 X_2 X_3 Y_0_NUDGED mlp
.options TEMP = 27
.options TNOM = 27
.tran 20ns 10665.6ns 0s
.end
