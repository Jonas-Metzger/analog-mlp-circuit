.title amp
Vin in 0 0V
Rin in mid 100Ohm
Bamp out 0 v={4 * (V(mid))}
Bdd mid 0 i={-0.25 * I(amp)}
Rout out 0 100Ohm
.options TEMP = 27
.options TNOM = 27
.dc Vin 0 1.95 0.01
.end
