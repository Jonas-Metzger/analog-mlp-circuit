.title Crossbar Circuit
.lib /root/miniforge3/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.subckt mlp NUDGED FREE X_0 X_1 X_2 Y_0_NUDGED Y_1_NUDGED
.subckt synapse WWL WBL RIN ROUT
Swrite_nfet MEM WBL WWL 0 switch
Ccap MEM ROUT 5.0pF capacitor
Mread_nfet ROUT MEM RIN RIN NMOSS l=5e-06 w=5e-06
.ends synapse

.subckt amplifier IN OUT
Bvcvs OUT 0 v={0 + 2 * (V(IN)-0)}
Bcccs INN 0 i={-0.5 * I(Bvcvs)}
Rmeas IN INN 0.001Ohm
Vdiou DIOU IN -0.25V
Ddiou DIOU 0 diode
.ends amplifier

.subckt optimizer1 WBL FREE NUDGED UPDATE NUDGED_OUTER
Bopamp OUT 0 v={V(WBL)*V(NUDGED_OUTER)/1.95}
Sstore OUT STORE NUDGED 0 switch
Cstore STORE 0 0.05pF capacitor
Sread STORE WBL UPDATE 0 switch
.ends optimizer1

.subckt optimizer100 WBL FREE NUDGED UPDATE NUDGED_OUTER
Bopamp OUT 0 v={V(WBL)*V(NUDGED_OUTER)/1.95}
Sstore OUT STORE NUDGED 0 switch
Cstore STORE 0 5.0pF capacitor
Sread STORE WBL UPDATE 0 switch
.ends optimizer100
Xweight_I0_H0 WWL_I0 WBL_IN_H0 X_0 IN_H0 synapse
Xweight_I1_H0 WWL_I1 WBL_IN_H0 X_1 IN_H0 synapse
Xweight_I2_H0 WWL_I2 WBL_IN_H0 X_2 IN_H0 synapse
Xact_H0 IN_H0 OUT_H0 amplifier
Xweight_J0_H0 WWL_J0 WBL_OUT_H0 OUT_H0 Y_0 synapse
Xweight_J1_H0 WWL_J1 WBL_OUT_H0 OUT_H0 Y_1 synapse
Xoptim_IN_H0 WBL_IN_H0 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H0 SET_IN_H0 WBL_IN_H0 SET 0 switch
SGND_IN_H0 IN_H0 0 SET 0 switch
Xoptim_OUT_H0 WBL_OUT_H0 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H0 SET_OUT_H0 WBL_OUT_H0 SET 0 switch
SGND_OUT_H0 OUT_H0 0 SET 0 switch
Xweight_I0_H1 WWL_I0 WBL_IN_H1 X_0 IN_H1 synapse
Xweight_I1_H1 WWL_I1 WBL_IN_H1 X_1 IN_H1 synapse
Xweight_I2_H1 WWL_I2 WBL_IN_H1 X_2 IN_H1 synapse
Xact_H1 IN_H1 OUT_H1 amplifier
Xweight_J0_H1 WWL_J0 WBL_OUT_H1 OUT_H1 Y_0 synapse
Xweight_J1_H1 WWL_J1 WBL_OUT_H1 OUT_H1 Y_1 synapse
Xoptim_IN_H1 WBL_IN_H1 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H1 SET_IN_H1 WBL_IN_H1 SET 0 switch
SGND_IN_H1 IN_H1 0 SET 0 switch
Xoptim_OUT_H1 WBL_OUT_H1 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H1 SET_OUT_H1 WBL_OUT_H1 SET 0 switch
SGND_OUT_H1 OUT_H1 0 SET 0 switch
Xweight_I0_H2 WWL_I0 WBL_IN_H2 X_0 IN_H2 synapse
Xweight_I1_H2 WWL_I1 WBL_IN_H2 X_1 IN_H2 synapse
Xweight_I2_H2 WWL_I2 WBL_IN_H2 X_2 IN_H2 synapse
Xact_H2 IN_H2 OUT_H2 amplifier
Xweight_J0_H2 WWL_J0 WBL_OUT_H2 OUT_H2 Y_0 synapse
Xweight_J1_H2 WWL_J1 WBL_OUT_H2 OUT_H2 Y_1 synapse
Xoptim_IN_H2 WBL_IN_H2 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H2 SET_IN_H2 WBL_IN_H2 SET 0 switch
SGND_IN_H2 IN_H2 0 SET 0 switch
Xoptim_OUT_H2 WBL_OUT_H2 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H2 SET_OUT_H2 WBL_OUT_H2 SET 0 switch
SGND_OUT_H2 OUT_H2 0 SET 0 switch
Xweight_I0_H3 WWL_I0 WBL_IN_H3 X_0 IN_H3 synapse
Xweight_I1_H3 WWL_I1 WBL_IN_H3 X_1 IN_H3 synapse
Xweight_I2_H3 WWL_I2 WBL_IN_H3 X_2 IN_H3 synapse
Xact_H3 IN_H3 OUT_H3 amplifier
Xweight_J0_H3 WWL_J0 WBL_OUT_H3 OUT_H3 Y_0 synapse
Xweight_J1_H3 WWL_J1 WBL_OUT_H3 OUT_H3 Y_1 synapse
Xoptim_IN_H3 WBL_IN_H3 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H3 SET_IN_H3 WBL_IN_H3 SET 0 switch
SGND_IN_H3 IN_H3 0 SET 0 switch
Xoptim_OUT_H3 WBL_OUT_H3 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H3 SET_OUT_H3 WBL_OUT_H3 SET 0 switch
SGND_OUT_H3 OUT_H3 0 SET 0 switch
Xweight_I0_H4 WWL_I0 WBL_IN_H4 X_0 IN_H4 synapse
Xweight_I1_H4 WWL_I1 WBL_IN_H4 X_1 IN_H4 synapse
Xweight_I2_H4 WWL_I2 WBL_IN_H4 X_2 IN_H4 synapse
Xact_H4 IN_H4 OUT_H4 amplifier
Xweight_J0_H4 WWL_J0 WBL_OUT_H4 OUT_H4 Y_0 synapse
Xweight_J1_H4 WWL_J1 WBL_OUT_H4 OUT_H4 Y_1 synapse
Xoptim_IN_H4 WBL_IN_H4 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H4 SET_IN_H4 WBL_IN_H4 SET 0 switch
SGND_IN_H4 IN_H4 0 SET 0 switch
Xoptim_OUT_H4 WBL_OUT_H4 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H4 SET_OUT_H4 WBL_OUT_H4 SET 0 switch
SGND_OUT_H4 OUT_H4 0 SET 0 switch
Xweight_I0_H5 WWL_I0 WBL_IN_H5 X_0 IN_H5 synapse
Xweight_I1_H5 WWL_I1 WBL_IN_H5 X_1 IN_H5 synapse
Xweight_I2_H5 WWL_I2 WBL_IN_H5 X_2 IN_H5 synapse
Xact_H5 IN_H5 OUT_H5 amplifier
Xweight_J0_H5 WWL_J0 WBL_OUT_H5 OUT_H5 Y_0 synapse
Xweight_J1_H5 WWL_J1 WBL_OUT_H5 OUT_H5 Y_1 synapse
Xoptim_IN_H5 WBL_IN_H5 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H5 SET_IN_H5 WBL_IN_H5 SET 0 switch
SGND_IN_H5 IN_H5 0 SET 0 switch
Xoptim_OUT_H5 WBL_OUT_H5 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H5 SET_OUT_H5 WBL_OUT_H5 SET 0 switch
SGND_OUT_H5 OUT_H5 0 SET 0 switch
Xweight_I0_H6 WWL_I0 WBL_IN_H6 X_0 IN_H6 synapse
Xweight_I1_H6 WWL_I1 WBL_IN_H6 X_1 IN_H6 synapse
Xweight_I2_H6 WWL_I2 WBL_IN_H6 X_2 IN_H6 synapse
Xact_H6 IN_H6 OUT_H6 amplifier
Xweight_J0_H6 WWL_J0 WBL_OUT_H6 OUT_H6 Y_0 synapse
Xweight_J1_H6 WWL_J1 WBL_OUT_H6 OUT_H6 Y_1 synapse
Xoptim_IN_H6 WBL_IN_H6 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H6 SET_IN_H6 WBL_IN_H6 SET 0 switch
SGND_IN_H6 IN_H6 0 SET 0 switch
Xoptim_OUT_H6 WBL_OUT_H6 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H6 SET_OUT_H6 WBL_OUT_H6 SET 0 switch
SGND_OUT_H6 OUT_H6 0 SET 0 switch
Xweight_I0_H7 WWL_I0 WBL_IN_H7 X_0 IN_H7 synapse
Xweight_I1_H7 WWL_I1 WBL_IN_H7 X_1 IN_H7 synapse
Xweight_I2_H7 WWL_I2 WBL_IN_H7 X_2 IN_H7 synapse
Xact_H7 IN_H7 OUT_H7 amplifier
Xweight_J0_H7 WWL_J0 WBL_OUT_H7 OUT_H7 Y_0 synapse
Xweight_J1_H7 WWL_J1 WBL_OUT_H7 OUT_H7 Y_1 synapse
Xoptim_IN_H7 WBL_IN_H7 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H7 SET_IN_H7 WBL_IN_H7 SET 0 switch
SGND_IN_H7 IN_H7 0 SET 0 switch
Xoptim_OUT_H7 WBL_OUT_H7 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H7 SET_OUT_H7 WBL_OUT_H7 SET 0 switch
SGND_OUT_H7 OUT_H7 0 SET 0 switch
Xweight_I0_H8 WWL_I0 WBL_IN_H8 X_0 IN_H8 synapse
Xweight_I1_H8 WWL_I1 WBL_IN_H8 X_1 IN_H8 synapse
Xweight_I2_H8 WWL_I2 WBL_IN_H8 X_2 IN_H8 synapse
Xact_H8 IN_H8 OUT_H8 amplifier
Xweight_J0_H8 WWL_J0 WBL_OUT_H8 OUT_H8 Y_0 synapse
Xweight_J1_H8 WWL_J1 WBL_OUT_H8 OUT_H8 Y_1 synapse
Xoptim_IN_H8 WBL_IN_H8 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H8 SET_IN_H8 WBL_IN_H8 SET 0 switch
SGND_IN_H8 IN_H8 0 SET 0 switch
Xoptim_OUT_H8 WBL_OUT_H8 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H8 SET_OUT_H8 WBL_OUT_H8 SET 0 switch
SGND_OUT_H8 OUT_H8 0 SET 0 switch
Xweight_I0_H9 WWL_I0 WBL_IN_H9 X_0 IN_H9 synapse
Xweight_I1_H9 WWL_I1 WBL_IN_H9 X_1 IN_H9 synapse
Xweight_I2_H9 WWL_I2 WBL_IN_H9 X_2 IN_H9 synapse
Xact_H9 IN_H9 OUT_H9 amplifier
Xweight_J0_H9 WWL_J0 WBL_OUT_H9 OUT_H9 Y_0 synapse
Xweight_J1_H9 WWL_J1 WBL_OUT_H9 OUT_H9 Y_1 synapse
Xoptim_IN_H9 WBL_IN_H9 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H9 SET_IN_H9 WBL_IN_H9 SET 0 switch
SGND_IN_H9 IN_H9 0 SET 0 switch
Xoptim_OUT_H9 WBL_OUT_H9 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H9 SET_OUT_H9 WBL_OUT_H9 SET 0 switch
SGND_OUT_H9 OUT_H9 0 SET 0 switch
Xweight_I0_H10 WWL_I0 WBL_IN_H10 X_0 IN_H10 synapse
Xweight_I1_H10 WWL_I1 WBL_IN_H10 X_1 IN_H10 synapse
Xweight_I2_H10 WWL_I2 WBL_IN_H10 X_2 IN_H10 synapse
Xact_H10 IN_H10 OUT_H10 amplifier
Xweight_J0_H10 WWL_J0 WBL_OUT_H10 OUT_H10 Y_0 synapse
Xweight_J1_H10 WWL_J1 WBL_OUT_H10 OUT_H10 Y_1 synapse
Xoptim_IN_H10 WBL_IN_H10 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H10 SET_IN_H10 WBL_IN_H10 SET 0 switch
SGND_IN_H10 IN_H10 0 SET 0 switch
Xoptim_OUT_H10 WBL_OUT_H10 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H10 SET_OUT_H10 WBL_OUT_H10 SET 0 switch
SGND_OUT_H10 OUT_H10 0 SET 0 switch
Xweight_I0_H11 WWL_I0 WBL_IN_H11 X_0 IN_H11 synapse
Xweight_I1_H11 WWL_I1 WBL_IN_H11 X_1 IN_H11 synapse
Xweight_I2_H11 WWL_I2 WBL_IN_H11 X_2 IN_H11 synapse
Xact_H11 IN_H11 OUT_H11 amplifier
Xweight_J0_H11 WWL_J0 WBL_OUT_H11 OUT_H11 Y_0 synapse
Xweight_J1_H11 WWL_J1 WBL_OUT_H11 OUT_H11 Y_1 synapse
Xoptim_IN_H11 WBL_IN_H11 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H11 SET_IN_H11 WBL_IN_H11 SET 0 switch
SGND_IN_H11 IN_H11 0 SET 0 switch
Xoptim_OUT_H11 WBL_OUT_H11 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H11 SET_OUT_H11 WBL_OUT_H11 SET 0 switch
SGND_OUT_H11 OUT_H11 0 SET 0 switch
Xweight_I0_H12 WWL_I0 WBL_IN_H12 X_0 IN_H12 synapse
Xweight_I1_H12 WWL_I1 WBL_IN_H12 X_1 IN_H12 synapse
Xweight_I2_H12 WWL_I2 WBL_IN_H12 X_2 IN_H12 synapse
Xact_H12 IN_H12 OUT_H12 amplifier
Xweight_J0_H12 WWL_J0 WBL_OUT_H12 OUT_H12 Y_0 synapse
Xweight_J1_H12 WWL_J1 WBL_OUT_H12 OUT_H12 Y_1 synapse
Xoptim_IN_H12 WBL_IN_H12 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H12 SET_IN_H12 WBL_IN_H12 SET 0 switch
SGND_IN_H12 IN_H12 0 SET 0 switch
Xoptim_OUT_H12 WBL_OUT_H12 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H12 SET_OUT_H12 WBL_OUT_H12 SET 0 switch
SGND_OUT_H12 OUT_H12 0 SET 0 switch
Xweight_I0_H13 WWL_I0 WBL_IN_H13 X_0 IN_H13 synapse
Xweight_I1_H13 WWL_I1 WBL_IN_H13 X_1 IN_H13 synapse
Xweight_I2_H13 WWL_I2 WBL_IN_H13 X_2 IN_H13 synapse
Xact_H13 IN_H13 OUT_H13 amplifier
Xweight_J0_H13 WWL_J0 WBL_OUT_H13 OUT_H13 Y_0 synapse
Xweight_J1_H13 WWL_J1 WBL_OUT_H13 OUT_H13 Y_1 synapse
Xoptim_IN_H13 WBL_IN_H13 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H13 SET_IN_H13 WBL_IN_H13 SET 0 switch
SGND_IN_H13 IN_H13 0 SET 0 switch
Xoptim_OUT_H13 WBL_OUT_H13 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H13 SET_OUT_H13 WBL_OUT_H13 SET 0 switch
SGND_OUT_H13 OUT_H13 0 SET 0 switch
Xweight_I0_H14 WWL_I0 WBL_IN_H14 X_0 IN_H14 synapse
Xweight_I1_H14 WWL_I1 WBL_IN_H14 X_1 IN_H14 synapse
Xweight_I2_H14 WWL_I2 WBL_IN_H14 X_2 IN_H14 synapse
Xact_H14 IN_H14 OUT_H14 amplifier
Xweight_J0_H14 WWL_J0 WBL_OUT_H14 OUT_H14 Y_0 synapse
Xweight_J1_H14 WWL_J1 WBL_OUT_H14 OUT_H14 Y_1 synapse
Xoptim_IN_H14 WBL_IN_H14 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H14 SET_IN_H14 WBL_IN_H14 SET 0 switch
SGND_IN_H14 IN_H14 0 SET 0 switch
Xoptim_OUT_H14 WBL_OUT_H14 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H14 SET_OUT_H14 WBL_OUT_H14 SET 0 switch
SGND_OUT_H14 OUT_H14 0 SET 0 switch
Xweight_I0_H15 WWL_I0 WBL_IN_H15 X_0 IN_H15 synapse
Xweight_I1_H15 WWL_I1 WBL_IN_H15 X_1 IN_H15 synapse
Xweight_I2_H15 WWL_I2 WBL_IN_H15 X_2 IN_H15 synapse
Xact_H15 IN_H15 OUT_H15 amplifier
Xweight_J0_H15 WWL_J0 WBL_OUT_H15 OUT_H15 Y_0 synapse
Xweight_J1_H15 WWL_J1 WBL_OUT_H15 OUT_H15 Y_1 synapse
Xoptim_IN_H15 WBL_IN_H15 FREE NUDGED UPDATE NUDGED_OUTER optimizer100
Sset_IN_H15 SET_IN_H15 WBL_IN_H15 SET 0 switch
SGND_IN_H15 IN_H15 0 SET 0 switch
Xoptim_OUT_H15 WBL_OUT_H15 FREE NUDGED UPDATE NUDGED_OUTER optimizer1
Sset_OUT_H15 SET_OUT_H15 WBL_OUT_H15 SET 0 switch
SGND_OUT_H15 OUT_H15 0 SET 0 switch
SY_0_NUDGED Y_0 Y_0_NUDGED NUDGED_OUTER 0 switch
SY_0_FREE Y_0 Y_0_FREE FREE 0 switch
CY_0_FREE Y_0_FREE 0 0.05pF capacitor
RY_0 Y_0 0 10kOhm
SY_1_NUDGED Y_1 Y_1_NUDGED NUDGED_OUTER 0 switch
SY_1_FREE Y_1 Y_1_FREE FREE 0 switch
CY_1_FREE Y_1_FREE 0 0.05pF capacitor
RY_1 Y_1 0 10kOhm
VSET_IN_H0 SET_IN_H0 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3237684667110443V 640000.0ns 0.3237684667110443V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.28780242800712585V 1520000.0ns 0.28780242800712585V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.3352009356021881V 2400000.0ns 0.3352009356021881V 2440000.0ns 0V)
VSET_OUT_H0 SET_OUT_H0 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.2941342294216156V 640000.0ns 0.2941342294216156V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.4893910884857178V 1520000.0ns 0.4893910884857178V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H1 SET_IN_H1 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.17695865035057068V 640000.0ns 0.17695865035057068V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.18991950154304504V 1520000.0ns 0.18991950154304504V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.47444629669189453V 2400000.0ns 0.47444629669189453V 2440000.0ns 0V)
VSET_OUT_H1 SET_OUT_H1 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.1070721372961998V 640000.0ns 0.1070721372961998V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.2985629141330719V 1520000.0ns 0.2985629141330719V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H2 SET_IN_H2 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.18539424240589142V 640000.0ns 0.18539424240589142V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.4309855103492737V 1520000.0ns 0.4309855103492737V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.33240142464637756V 2400000.0ns 0.33240142464637756V 2440000.0ns 0V)
VSET_OUT_H2 SET_OUT_H2 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3552550673484802V 640000.0ns 0.3552550673484802V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.19294896721839905V 1520000.0ns 0.19294896721839905V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H3 SET_IN_H3 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.24866893887519836V 640000.0ns 0.24866893887519836V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.3644316792488098V 1520000.0ns 0.3644316792488098V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.154496431350708V 2400000.0ns 0.154496431350708V 2440000.0ns 0V)
VSET_OUT_H3 SET_OUT_H3 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.18904300034046173V 640000.0ns 0.18904300034046173V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.4340851306915283V 1520000.0ns 0.4340851306915283V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H4 SET_IN_H4 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.36711385846138V 640000.0ns 0.36711385846138V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.13436710834503174V 1520000.0ns 0.13436710834503174V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.18623051047325134V 2400000.0ns 0.18623051047325134V 2440000.0ns 0V)
VSET_OUT_H4 SET_OUT_H4 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.17669212818145752V 640000.0ns 0.17669212818145752V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.46766600012779236V 1520000.0ns 0.46766600012779236V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H5 SET_IN_H5 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3603936433792114V 640000.0ns 0.3603936433792114V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.31234630942344666V 1520000.0ns 0.31234630942344666V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.20562931895256042V 2400000.0ns 0.20562931895256042V 2440000.0ns 0V)
VSET_OUT_H5 SET_OUT_H5 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.282827764749527V 640000.0ns 0.282827764749527V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.20167246460914612V 1520000.0ns 0.20167246460914612V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H6 SET_IN_H6 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.268454372882843V 640000.0ns 0.268454372882843V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.41979044675827026V 1520000.0ns 0.41979044675827026V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.3936837613582611V 2400000.0ns 0.3936837613582611V 2440000.0ns 0V)
VSET_OUT_H6 SET_OUT_H6 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.39986422657966614V 640000.0ns 0.39986422657966614V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.1662781983613968V 1520000.0ns 0.1662781983613968V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H7 SET_IN_H7 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3497702479362488V 640000.0ns 0.3497702479362488V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.35625243186950684V 1520000.0ns 0.35625243186950684V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.20707571506500244V 2400000.0ns 0.20707571506500244V 2440000.0ns 0V)
VSET_OUT_H7 SET_OUT_H7 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.30827999114990234V 640000.0ns 0.30827999114990234V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.44093620777130127V 1520000.0ns 0.44093620777130127V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H8 SET_IN_H8 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.49417197704315186V 640000.0ns 0.49417197704315186V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.16059112548828125V 1520000.0ns 0.16059112548828125V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.17716260254383087V 2400000.0ns 0.17716260254383087V 2440000.0ns 0V)
VSET_OUT_H8 SET_OUT_H8 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3837760090827942V 640000.0ns 0.3837760090827942V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.3614835739135742V 1520000.0ns 0.3614835739135742V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H9 SET_IN_H9 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.2293718457221985V 640000.0ns 0.2293718457221985V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.2944580018520355V 1520000.0ns 0.2944580018520355V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.39146584272384644V 2400000.0ns 0.39146584272384644V 2440000.0ns 0V)
VSET_OUT_H9 SET_OUT_H9 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.46183472871780396V 640000.0ns 0.46183472871780396V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.38461968302726746V 1520000.0ns 0.38461968302726746V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H10 SET_IN_H10 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.37664541602134705V 640000.0ns 0.37664541602134705V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.12331042438745499V 1520000.0ns 0.12331042438745499V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.19100043177604675V 2400000.0ns 0.19100043177604675V 2440000.0ns 0V)
VSET_OUT_H10 SET_OUT_H10 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3277418911457062V 640000.0ns 0.3277418911457062V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.3207624852657318V 1520000.0ns 0.3207624852657318V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H11 SET_IN_H11 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.17984595894813538V 640000.0ns 0.17984595894813538V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.2194565236568451V 1520000.0ns 0.2194565236568451V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.2143402397632599V 2400000.0ns 0.2143402397632599V 2440000.0ns 0V)
VSET_OUT_H11 SET_OUT_H11 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.34952303767204285V 640000.0ns 0.34952303767204285V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.4432114064693451V 1520000.0ns 0.4432114064693451V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H12 SET_IN_H12 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.2933448255062103V 640000.0ns 0.2933448255062103V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.11042072623968124V 1520000.0ns 0.11042072623968124V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.49986961483955383V 2400000.0ns 0.49986961483955383V 2440000.0ns 0V)
VSET_OUT_H12 SET_OUT_H12 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.4447947144508362V 640000.0ns 0.4447947144508362V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.12481585144996643V 1520000.0ns 0.12481585144996643V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H13 SET_IN_H13 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3627299666404724V 640000.0ns 0.3627299666404724V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.10622155666351318V 1520000.0ns 0.10622155666351318V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.12430758774280548V 2400000.0ns 0.12430758774280548V 2440000.0ns 0V)
VSET_OUT_H13 SET_OUT_H13 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.2213345319032669V 640000.0ns 0.2213345319032669V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.13766613602638245V 1520000.0ns 0.13766613602638245V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H14 SET_IN_H14 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.20897206664085388V 640000.0ns 0.20897206664085388V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.46652302145957947V 1520000.0ns 0.46652302145957947V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.4699414372444153V 2400000.0ns 0.4699414372444153V 2440000.0ns 0V)
VSET_OUT_H14 SET_OUT_H14 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.4986300766468048V 640000.0ns 0.4986300766468048V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.4820975363254547V 1520000.0ns 0.4820975363254547V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET_IN_H15 SET_IN_H15 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.15766611695289612V 640000.0ns 0.15766611695289612V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.20440998673439026V 1520000.0ns 0.20440998673439026V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0.3871707320213318V 2400000.0ns 0.3871707320213318V 2440000.0ns 0V)
VSET_OUT_H15 SET_OUT_H15 0 PWL(0ns 0V 200000.0ns 0V 240000.0ns 0.3147434890270233V 640000.0ns 0.3147434890270233V 680000.0ns 0V 1080000.0ns 0V 1120000.0ns 0.4686463475227356V 1520000.0ns 0.4686463475227356V 1560000.0ns 0V 1960000.0ns 0V 2000000.0ns 0V 2400000.0ns 0V 2440000.0ns 0V)
VSET SET 0 PWL(0ns 1.95V 3080000.0ns 1.95V 3120000.0ns 0V)
VNUDGED NUDGED 0 PWL(0ns 0V 3960000.0ns 0V 7800000.0ns 0V 7840000.0ns 0V 8240000.0ns 0V 8280000.0ns 0V 9080000.0ns 0V 9120000.0ns 1.95V 9520000.0ns 1.95V 9560000.0ns 0V 10360000.0ns 0V 10400000.0ns 0V 10800000.0ns 0V 10840000.0ns 0V 11640000.0ns 0V 11680000.0ns 0V 12080000.0ns 0V 12120000.0ns 0V 12920000.0ns 0V 12960000.0ns 1.95V 13360000.0ns 1.95V 13400000.0ns 0V 14200000.0ns 0V 14240000.0ns 0V 14640000.0ns 0V 14680000.0ns 0V 15480000.0ns 0V 15520000.0ns 0V 15920000.0ns 0V 15960000.0ns 0V 16760000.0ns 0V 16800000.0ns 1.95V 17200000.0ns 1.95V 17240000.0ns 0V 18040000.0ns 0V 18080000.0ns 0V 18480000.0ns 0V 18520000.0ns 0V 19320000.0ns 0V 19360000.0ns 0V 19760000.0ns 0V 19800000.0ns 0V 20600000.0ns 0V 20640000.0ns 1.95V 21040000.0ns 1.95V 21080000.0ns 0V 21880000.0ns 0V 21920000.0ns 0V 22320000.0ns 0V 22360000.0ns 0V 23160000.0ns 0V 23200000.0ns 0V 23600000.0ns 0V 23640000.0ns 0V 24440000.0ns 0V 24480000.0ns 1.95V 24880000.0ns 1.95V 24920000.0ns 0V 25720000.0ns 0V 25760000.0ns 0V 26160000.0ns 0V 26200000.0ns 0V 27000000.0ns 0V 27040000.0ns 0V 27440000.0ns 0V 27480000.0ns 0V 28280000.0ns 0V 28320000.0ns 1.95V 28720000.0ns 1.95V 28760000.0ns 0V 29560000.0ns 0V 29600000.0ns 0V 30000000.0ns 0V 30040000.0ns 0V 30840000.0ns 0V 30880000.0ns 0V 31280000.0ns 0V 31320000.0ns 0V 32120000.0ns 0V 32160000.0ns 1.95V 32560000.0ns 1.95V 32600000.0ns 0V 33400000.0ns 0V 33440000.0ns 0V 33840000.0ns 0V 33880000.0ns 0V 34680000.0ns 0V 34720000.0ns 0V 35120000.0ns 0V 35160000.0ns 0V 35960000.0ns 0V 36000000.0ns 1.95V 36400000.0ns 1.95V 36440000.0ns 0V 37240000.0ns 0V 37280000.0ns 0V 37680000.0ns 0V 37720000.0ns 0V 38520000.0ns 0V 38560000.0ns 0V 38960000.0ns 0V 39000000.0ns 0V 39800000.0ns 0V 39840000.0ns 1.95V 40240000.0ns 1.95V 40280000.0ns 0V 41080000.0ns 0V 41120000.0ns 0V 41520000.0ns 0V 41560000.0ns 0V 42360000.0ns 0V 42400000.0ns 0V 42800000.0ns 0V 42840000.0ns 0V 43640000.0ns 0V 43680000.0ns 1.95V 44080000.0ns 1.95V 44120000.0ns 0V 44920000.0ns 0V 44960000.0ns 0V 45360000.0ns 0V 45400000.0ns 0V 46200000.0ns 0V 46240000.0ns 0V 46640000.0ns 0V 46680000.0ns 0V 47480000.0ns 0V 47520000.0ns 1.95V 47920000.0ns 1.95V 47960000.0ns 0V 48760000.0ns 0V 48800000.0ns 0V 49200000.0ns 0V 49240000.0ns 0V 50040000.0ns 0V 50080000.0ns 0V 50480000.0ns 0V 50520000.0ns 0V 51320000.0ns 0V 51360000.0ns 1.95V 51760000.0ns 1.95V 51800000.0ns 0V 52600000.0ns 0V 52640000.0ns 0V 53040000.0ns 0V 53080000.0ns 0V 53880000.0ns 0V 53920000.0ns 0V 54320000.0ns 0V 54360000.0ns 0V 55160000.0ns 0V 55200000.0ns 1.95V 55600000.0ns 1.95V 55640000.0ns 0V 56440000.0ns 0V 56480000.0ns 0V 56880000.0ns 0V 56920000.0ns 0V 57720000.0ns 0V 57760000.0ns 0V 58160000.0ns 0V 58200000.0ns 0V 59000000.0ns 0V 59040000.0ns 1.95V 59440000.0ns 1.95V 59480000.0ns 0V 60280000.0ns 0V 60320000.0ns 0V 60720000.0ns 0V 60760000.0ns 0V 61560000.0ns 0V 61600000.0ns 0V 62000000.0ns 0V 62040000.0ns 0V 62840000.0ns 0V 62880000.0ns 1.95V 63280000.0ns 1.95V 63320000.0ns 0V 64120000.0ns 0V 64160000.0ns 0V 64560000.0ns 0V 64600000.0ns 0V 65400000.0ns 0V 65440000.0ns 0V 65840000.0ns 0V 65880000.0ns 0V 66680000.0ns 0V 66720000.0ns 1.95V 67120000.0ns 1.95V 67160000.0ns 0V 67960000.0ns 0V 68000000.0ns 0V 68400000.0ns 0V 68440000.0ns 0V 69240000.0ns 0V 69280000.0ns 0V 69680000.0ns 0V 69720000.0ns 0V 70520000.0ns 0V 70560000.0ns 1.95V 70960000.0ns 1.95V 71000000.0ns 0V 71800000.0ns 0V 71840000.0ns 0V 72240000.0ns 0V 72280000.0ns 0V 73080000.0ns 0V 73120000.0ns 0V 73520000.0ns 0V 73560000.0ns 0V 74360000.0ns 0V 74400000.0ns 1.95V 74800000.0ns 1.95V 74840000.0ns 0V 75640000.0ns 0V 75680000.0ns 0V 76080000.0ns 0V 76120000.0ns 0V 76920000.0ns 0V 76960000.0ns 0V 77360000.0ns 0V 77400000.0ns 0V 78200000.0ns 0V 78240000.0ns 1.95V 78640000.0ns 1.95V 78680000.0ns 0V 79480000.0ns 0V 79520000.0ns 0V 79920000.0ns 0V 79960000.0ns 0V 80760000.0ns 0V 80800000.0ns 0V 81200000.0ns 0V 81240000.0ns 0V 82040000.0ns 0V 82080000.0ns 1.95V 82480000.0ns 1.95V 82520000.0ns 0V 83320000.0ns 0V 83360000.0ns 0V 83760000.0ns 0V 83800000.0ns 0V 84600000.0ns 0V 84640000.0ns 0V 85040000.0ns 0V 85080000.0ns 0V 85880000.0ns 0V 85920000.0ns 1.95V 86320000.0ns 1.95V 86360000.0ns 0V 87160000.0ns 0V 87200000.0ns 0V 87600000.0ns 0V 87640000.0ns 0V 88440000.0ns 0V 88480000.0ns 0V 88880000.0ns 0V 88920000.0ns 0V 89720000.0ns 0V 89760000.0ns 1.95V 90160000.0ns 1.95V 90200000.0ns 0V 91000000.0ns 0V 91040000.0ns 0V 91440000.0ns 0V 91480000.0ns 0V 92280000.0ns 0V 92320000.0ns 0V 92720000.0ns 0V 92760000.0ns 0V 93560000.0ns 0V 93600000.0ns 1.95V 94000000.0ns 1.95V 94040000.0ns 0V 94840000.0ns 0V 94880000.0ns 0V 95280000.0ns 0V 95320000.0ns 0V 96120000.0ns 0V 96160000.0ns 0V 96560000.0ns 0V 96600000.0ns 0V 97400000.0ns 0V 97440000.0ns 1.95V 97840000.0ns 1.95V 97880000.0ns 0V 98680000.0ns 0V 98720000.0ns 0V 99120000.0ns 0V 99160000.0ns 0V 99960000.0ns 0V 100000000.0ns 0V 100400000.0ns 0V 100440000.0ns 0V 101240000.0ns 0V 101280000.0ns 1.95V 101680000.0ns 1.95V 101720000.0ns 0V 102520000.0ns 0V 102560000.0ns 0V 102960000.0ns 0V 103000000.0ns 0V 103800000.0ns 0V 103840000.0ns 0V 104240000.0ns 0V 104280000.0ns 0V 105080000.0ns 0V 105120000.0ns 1.95V 105520000.0ns 1.95V 105560000.0ns 0V 106360000.0ns 0V 106400000.0ns 0V 106800000.0ns 0V 106840000.0ns 0V 107640000.0ns 0V 107680000.0ns 0V 108080000.0ns 0V 108120000.0ns 0V 108920000.0ns 0V 108960000.0ns 1.95V 109360000.0ns 1.95V 109400000.0ns 0V 110200000.0ns 0V 110240000.0ns 0V 110640000.0ns 0V 110680000.0ns 0V 111480000.0ns 0V 111520000.0ns 0V 111920000.0ns 0V 111960000.0ns 0V 112760000.0ns 0V 112800000.0ns 1.95V 113200000.0ns 1.95V 113240000.0ns 0V 114040000.0ns 0V 114080000.0ns 0V 114480000.0ns 0V 114520000.0ns 0V 115320000.0ns 0V 115360000.0ns 0V 115760000.0ns 0V 115800000.0ns 0V 116600000.0ns 0V 116640000.0ns 1.95V 117040000.0ns 1.95V 117080000.0ns 0V 117880000.0ns 0V 117920000.0ns 0V 118320000.0ns 0V 118360000.0ns 0V 119160000.0ns 0V 119200000.0ns 0V 119600000.0ns 0V 119640000.0ns 0V 120440000.0ns 0V 120480000.0ns 1.95V 120880000.0ns 1.95V 120920000.0ns 0V 121720000.0ns 0V 121760000.0ns 0V 122160000.0ns 0V 122200000.0ns 0V 123000000.0ns 0V 123040000.0ns 0V 123440000.0ns 0V 123480000.0ns 0V 124280000.0ns 0V 124320000.0ns 1.95V 124720000.0ns 1.95V 124760000.0ns 0V 125560000.0ns 0V 125600000.0ns 0V 126000000.0ns 0V 126040000.0ns 0V 126840000.0ns 0V 126880000.0ns 0V 127280000.0ns 0V 127320000.0ns 0V 128120000.0ns 0V 128160000.0ns 1.95V 128560000.0ns 1.95V 128600000.0ns 0V 129400000.0ns 0V 129440000.0ns 0V 129840000.0ns 0V 129880000.0ns 0V 130680000.0ns 0V 130720000.0ns 0V 131120000.0ns 0V 131160000.0ns 0V 131960000.0ns 0V 132000000.0ns 1.95V 132400000.0ns 1.95V 132440000.0ns 0V 133240000.0ns 0V 133280000.0ns 0V 133680000.0ns 0V 133720000.0ns 0V 134520000.0ns 0V 134560000.0ns 0V 134960000.0ns 0V 135000000.0ns 0V 135800000.0ns 0V 135840000.0ns 1.95V 136240000.0ns 1.95V 136280000.0ns 0V 137080000.0ns 0V 137120000.0ns 0V 137520000.0ns 0V 137560000.0ns 0V 138360000.0ns 0V 138400000.0ns 0V 138800000.0ns 0V 138840000.0ns 0V 139640000.0ns 0V 139680000.0ns 1.95V 140080000.0ns 1.95V 140120000.0ns 0V 140920000.0ns 0V 140960000.0ns 0V 141360000.0ns 0V 141400000.0ns 0V 142200000.0ns 0V 142240000.0ns 0V 142640000.0ns 0V 142680000.0ns 0V 143480000.0ns 0V 143520000.0ns 1.95V 143920000.0ns 1.95V 143960000.0ns 0V 144760000.0ns 0V 144800000.0ns 0V 145200000.0ns 0V 145240000.0ns 0V 146040000.0ns 0V 146080000.0ns 0V 146480000.0ns 0V 146520000.0ns 0V 147320000.0ns 0V 147360000.0ns 1.95V 147760000.0ns 1.95V 147800000.0ns 0V 148600000.0ns 0V 148640000.0ns 0V 149040000.0ns 0V 149080000.0ns 0V 149880000.0ns 0V 149920000.0ns 0V 150320000.0ns 0V 150360000.0ns 0V 151160000.0ns 0V 151200000.0ns 1.95V 151600000.0ns 1.95V 151640000.0ns 0V 152440000.0ns 0V 152480000.0ns 0V 152880000.0ns 0V 152920000.0ns 0V 153720000.0ns 0V 153760000.0ns 0V 154160000.0ns 0V 154200000.0ns 0V 155000000.0ns 0V 155040000.0ns 1.95V 155440000.0ns 1.95V 155480000.0ns 0V 156280000.0ns 0V 156320000.0ns 0V 156720000.0ns 0V 156760000.0ns 0V 157560000.0ns 0V 157600000.0ns 0V 158000000.0ns 0V 158040000.0ns 0V 158840000.0ns 0V 158880000.0ns 1.95V 159280000.0ns 1.95V 159320000.0ns 0V 160120000.0ns 0V 160160000.0ns 0V 160560000.0ns 0V 160600000.0ns 0V 161400000.0ns 0V 161440000.0ns 0V 161840000.0ns 0V 161880000.0ns 0V 162680000.0ns 0V 162720000.0ns 1.95V 163120000.0ns 1.95V 163160000.0ns 0V 163960000.0ns 0V 164000000.0ns 0V 164400000.0ns 0V 164440000.0ns 0V 165240000.0ns 0V 165280000.0ns 0V 165680000.0ns 0V 165720000.0ns 0V 166520000.0ns 0V 166560000.0ns 1.95V 166960000.0ns 1.95V 167000000.0ns 0V 167800000.0ns 0V 167840000.0ns 0V 168240000.0ns 0V 168280000.0ns 0V 169080000.0ns 0V 169120000.0ns 0V 169520000.0ns 0V 169560000.0ns 0V 170360000.0ns 0V 170400000.0ns 1.95V 170800000.0ns 1.95V 170840000.0ns 0V 171640000.0ns 0V 171680000.0ns 0V 172080000.0ns 0V 172120000.0ns 0V 172920000.0ns 0V 172960000.0ns 0V 173360000.0ns 0V 173400000.0ns 0V 174200000.0ns 0V 174240000.0ns 1.95V 174640000.0ns 1.95V 174680000.0ns 0V 175480000.0ns 0V 175520000.0ns 0V 175920000.0ns 0V 175960000.0ns 0V 176760000.0ns 0V 176800000.0ns 0V 177200000.0ns 0V 177240000.0ns 0V 178040000.0ns 0V 178080000.0ns 1.95V 178480000.0ns 1.95V 178520000.0ns 0V 179320000.0ns 0V 179360000.0ns 0V 179760000.0ns 0V 179800000.0ns 0V 180600000.0ns 0V 180640000.0ns 0V 181040000.0ns 0V 181080000.0ns 0V 181880000.0ns 0V 181920000.0ns 1.95V 182320000.0ns 1.95V 182360000.0ns 0V 183160000.0ns 0V 183200000.0ns 0V 183600000.0ns 0V 183640000.0ns 0V 184440000.0ns 0V 184480000.0ns 0V 184880000.0ns 0V 184920000.0ns 0V 185720000.0ns 0V 185760000.0ns 1.95V 186160000.0ns 1.95V 186200000.0ns 0V 187000000.0ns 0V 187040000.0ns 0V 187440000.0ns 0V 187480000.0ns 0V 188280000.0ns 0V 188320000.0ns 0V 188720000.0ns 0V 188760000.0ns 0V 189560000.0ns 0V 189600000.0ns 1.95V 190000000.0ns 1.95V 190040000.0ns 0V 190840000.0ns 0V 190880000.0ns 0V 191280000.0ns 0V 191320000.0ns 0V 192120000.0ns 0V 192160000.0ns 0V 192560000.0ns 0V 192600000.0ns 0V 193400000.0ns 0V 193440000.0ns 1.95V 193840000.0ns 1.95V 193880000.0ns 0V 194680000.0ns 0V 194720000.0ns 0V 195120000.0ns 0V 195160000.0ns 0V 195960000.0ns 0V 196000000.0ns 0V 196400000.0ns 0V 196440000.0ns 0V 197240000.0ns 0V 197280000.0ns 1.95V 197680000.0ns 1.95V 197720000.0ns 0V 198520000.0ns 0V 198560000.0ns 0V 198960000.0ns 0V 199000000.0ns 0V 199800000.0ns 0V 199840000.0ns 0V 200240000.0ns 0V 200280000.0ns 0V 201080000.0ns 0V 201120000.0ns 1.95V 201520000.0ns 1.95V 201560000.0ns 0V 202360000.0ns 0V 202400000.0ns 0V 202800000.0ns 0V 202840000.0ns 0V 203640000.0ns 0V 203680000.0ns 0V 204080000.0ns 0V 204120000.0ns 0V 204920000.0ns 0V 204960000.0ns 1.95V 205360000.0ns 1.95V 205400000.0ns 0V 206200000.0ns 0V 206240000.0ns 0V 206640000.0ns 0V 206680000.0ns 0V 207480000.0ns 0V 207520000.0ns 0V 207920000.0ns 0V 207960000.0ns 0V 208760000.0ns 0V 208800000.0ns 1.95V 209200000.0ns 1.95V 209240000.0ns 0V 210040000.0ns 0V 210080000.0ns 0V 210480000.0ns 0V 210520000.0ns 0V 211320000.0ns 0V 211360000.0ns 0V 211760000.0ns 0V 211800000.0ns 0V 212600000.0ns 0V 212640000.0ns 1.95V 213040000.0ns 1.95V 213080000.0ns 0V 213880000.0ns 0V 213920000.0ns 0V 214320000.0ns 0V 214360000.0ns 0V 215160000.0ns 0V 215200000.0ns 0V 215600000.0ns 0V 215640000.0ns 0V 216440000.0ns 0V 216480000.0ns 1.95V 216880000.0ns 1.95V 216920000.0ns 0V 217720000.0ns 0V 217760000.0ns 0V 218160000.0ns 0V 218200000.0ns 0V 219000000.0ns 0V 219040000.0ns 0V 219440000.0ns 0V 219480000.0ns 0V 220280000.0ns 0V 220320000.0ns 1.95V 220720000.0ns 1.95V 220760000.0ns 0V 221560000.0ns 0V 221600000.0ns 0V 222000000.0ns 0V 222040000.0ns 0V 222840000.0ns 0V 222880000.0ns 0V 223280000.0ns 0V 223320000.0ns 0V 224120000.0ns 0V 224160000.0ns 1.95V 224560000.0ns 1.95V 224600000.0ns 0V 225400000.0ns 0V 225440000.0ns 0V 225840000.0ns 0V 225880000.0ns 0V 226680000.0ns 0V 226720000.0ns 0V 227120000.0ns 0V 227160000.0ns 0V 227960000.0ns 0V 228000000.0ns 1.95V 228400000.0ns 1.95V 228440000.0ns 0V 229240000.0ns 0V 229280000.0ns 0V 229680000.0ns 0V 229720000.0ns 0V 230520000.0ns 0V 230560000.0ns 0V 230960000.0ns 0V 231000000.0ns 0V 231800000.0ns 0V 231840000.0ns 1.95V 232240000.0ns 1.95V 232280000.0ns 0V 233080000.0ns 0V 233120000.0ns 0V 233520000.0ns 0V 233560000.0ns 0V 234360000.0ns 0V 234400000.0ns 0V 234800000.0ns 0V 234840000.0ns 0V 235640000.0ns 0V 235680000.0ns 1.95V 236080000.0ns 1.95V 236120000.0ns 0V 236920000.0ns 0V 236960000.0ns 0V 237360000.0ns 0V 237400000.0ns 0V 238200000.0ns 0V 238240000.0ns 0V 238640000.0ns 0V 238680000.0ns 0V 239480000.0ns 0V 239520000.0ns 1.95V 239920000.0ns 1.95V 239960000.0ns 0V 240760000.0ns 0V 240800000.0ns 0V 241200000.0ns 0V 241240000.0ns 0V 242040000.0ns 0V 242080000.0ns 0V 242480000.0ns 0V 242520000.0ns 0V 243320000.0ns 0V 243360000.0ns 1.95V 243760000.0ns 1.95V 243800000.0ns 0V 244600000.0ns 0V 244640000.0ns 0V 245040000.0ns 0V 245080000.0ns 0V 245880000.0ns 0V 245920000.0ns 0V 246320000.0ns 0V 246360000.0ns 0V 247160000.0ns 0V 247200000.0ns 1.95V 247600000.0ns 1.95V 247640000.0ns 0V 248440000.0ns 0V 248480000.0ns 0V 248880000.0ns 0V 248920000.0ns 0V 249720000.0ns 0V 249760000.0ns 0V 250160000.0ns 0V 250200000.0ns 0V 251000000.0ns 0V 251040000.0ns 1.95V 251440000.0ns 1.95V 251480000.0ns 0V 252280000.0ns 0V 252320000.0ns 0V 252720000.0ns 0V 252760000.0ns 0V 253560000.0ns 0V 253600000.0ns 0V 254000000.0ns 0V 254040000.0ns 0V 254840000.0ns 0V 254880000.0ns 1.95V 255280000.0ns 1.95V 255320000.0ns 0V 256120000.0ns 0V 256160000.0ns 0V 256560000.0ns 0V 256600000.0ns 0V 257400000.0ns 0V 257440000.0ns 0V 257840000.0ns 0V 257880000.0ns 0V 258680000.0ns 0V 258720000.0ns 1.95V 259120000.0ns 1.95V 259160000.0ns 0V 259960000.0ns 0V 260000000.0ns 0V 260400000.0ns 0V 260440000.0ns 0V 261240000.0ns 0V 261280000.0ns 0V 261680000.0ns 0V 261720000.0ns 0V 262520000.0ns 0V 262560000.0ns 1.95V 262960000.0ns 1.95V 263000000.0ns 0V 263800000.0ns 0V 263840000.0ns 0V 264240000.0ns 0V 264280000.0ns 0V 265080000.0ns 0V 265120000.0ns 0V 265520000.0ns 0V 265560000.0ns 0V 266360000.0ns 0V 266400000.0ns 1.95V 266800000.0ns 1.95V 266840000.0ns 0V 267640000.0ns 0V 267680000.0ns 0V 268080000.0ns 0V 268120000.0ns 0V 268920000.0ns 0V 268960000.0ns 0V 269360000.0ns 0V 269400000.0ns 0V 270200000.0ns 0V 270240000.0ns 1.95V 270640000.0ns 1.95V 270680000.0ns 0V 271480000.0ns 0V 271520000.0ns 0V 271920000.0ns 0V 271960000.0ns 0V 272760000.0ns 0V 272800000.0ns 0V 273200000.0ns 0V 273240000.0ns 0V 274040000.0ns 0V 274080000.0ns 1.95V 274480000.0ns 1.95V 274520000.0ns 0V 275320000.0ns 0V 275360000.0ns 0V 275760000.0ns 0V 275800000.0ns 0V 276600000.0ns 0V 276640000.0ns 0V 277040000.0ns 0V 277080000.0ns 0V 277880000.0ns 0V 277920000.0ns 1.95V 278320000.0ns 1.95V 278360000.0ns 0V 279160000.0ns 0V 279200000.0ns 0V 279600000.0ns 0V 279640000.0ns 0V 280440000.0ns 0V 280480000.0ns 0V 280880000.0ns 0V 280920000.0ns 0V 281720000.0ns 0V 281760000.0ns 1.95V 282160000.0ns 1.95V 282200000.0ns 0V 283000000.0ns 0V 283040000.0ns 0V 283440000.0ns 0V 283480000.0ns 0V 284280000.0ns 0V 284320000.0ns 0V 284720000.0ns 0V 284760000.0ns 0V 285560000.0ns 0V 285600000.0ns 1.95V 286000000.0ns 1.95V 286040000.0ns 0V 286840000.0ns 0V 286880000.0ns 0V 287280000.0ns 0V 287320000.0ns 0V 288120000.0ns 0V 288160000.0ns 0V 288560000.0ns 0V 288600000.0ns 0V 289400000.0ns 0V 289440000.0ns 1.95V 289840000.0ns 1.95V 289880000.0ns 0V 290680000.0ns 0V 290720000.0ns 0V 291120000.0ns 0V 291160000.0ns 0V 291960000.0ns 0V 292000000.0ns 0V 292400000.0ns 0V 292440000.0ns 0V 293240000.0ns 0V 293280000.0ns 1.95V 293680000.0ns 1.95V 293720000.0ns 0V 294520000.0ns 0V 294560000.0ns 0V 294960000.0ns 0V 295000000.0ns 0V 295800000.0ns 0V 295840000.0ns 0V 296240000.0ns 0V 296280000.0ns 0V 297080000.0ns 0V 297120000.0ns 1.95V 297520000.0ns 1.95V 297560000.0ns 0V 298360000.0ns 0V 298400000.0ns 0V 298800000.0ns 0V 298840000.0ns 0V 299640000.0ns 0V 299680000.0ns 0V 300080000.0ns 0V 300120000.0ns 0V 300920000.0ns 0V 300960000.0ns 1.95V 301360000.0ns 1.95V 301400000.0ns 0V 302200000.0ns 0V 302240000.0ns 0V 302640000.0ns 0V 302680000.0ns 0V 303480000.0ns 0V 303520000.0ns 0V 303920000.0ns 0V 303960000.0ns 0V 304760000.0ns 0V 304800000.0ns 1.95V 305200000.0ns 1.95V 305240000.0ns 0V 306040000.0ns 0V 306080000.0ns 0V 306480000.0ns 0V 306520000.0ns 0V 307320000.0ns 0V 307360000.0ns 0V 307760000.0ns 0V 307800000.0ns 0V 308600000.0ns 0V 308640000.0ns 1.95V 309040000.0ns 1.95V 309080000.0ns 0V 309880000.0ns 0V 309920000.0ns 0V 310320000.0ns 0V 310360000.0ns 0V 311160000.0ns 0V 311200000.0ns 0V 311600000.0ns 0V 311640000.0ns 0V 312440000.0ns 0V 312480000.0ns 1.95V 312880000.0ns 1.95V 312920000.0ns 0V 313720000.0ns 0V 313760000.0ns 0V 314160000.0ns 0V 314200000.0ns 0V 315000000.0ns 0V 315040000.0ns 0V 315440000.0ns 0V 315480000.0ns 0V 316280000.0ns 0V 316320000.0ns 1.95V 316720000.0ns 1.95V 316760000.0ns 0V 317560000.0ns 0V 317600000.0ns 0V 318000000.0ns 0V 318040000.0ns 0V 318840000.0ns 0V 318880000.0ns 0V 319280000.0ns 0V 319320000.0ns 0V 320120000.0ns 0V 320160000.0ns 1.95V 320560000.0ns 1.95V 320600000.0ns 0V 321400000.0ns 0V 321440000.0ns 0V 321840000.0ns 0V 321880000.0ns 0V 322680000.0ns 0V 322720000.0ns 0V 323120000.0ns 0V 323160000.0ns 0V 323960000.0ns 0V 324000000.0ns 1.95V 324400000.0ns 1.95V 324440000.0ns 0V 325240000.0ns 0V 325280000.0ns 0V 325680000.0ns 0V 325720000.0ns 0V 326520000.0ns 0V 326560000.0ns 0V 326960000.0ns 0V 327000000.0ns 0V 327800000.0ns 0V 327840000.0ns 1.95V 328240000.0ns 1.95V 328280000.0ns 0V 329080000.0ns 0V 329120000.0ns 0V 329520000.0ns 0V 329560000.0ns 0V 330360000.0ns 0V 330400000.0ns 0V 330800000.0ns 0V 330840000.0ns 0V 331640000.0ns 0V 331680000.0ns 1.95V 332080000.0ns 1.95V 332120000.0ns 0V 332920000.0ns 0V 332960000.0ns 0V 333360000.0ns 0V 333400000.0ns 0V 334200000.0ns 0V 334240000.0ns 0V 334640000.0ns 0V 334680000.0ns 0V 335480000.0ns 0V 335520000.0ns 1.95V 335920000.0ns 1.95V 335960000.0ns 0V 336760000.0ns 0V 336800000.0ns 0V 337200000.0ns 0V 337240000.0ns 0V 338040000.0ns 0V 338080000.0ns 0V 338480000.0ns 0V 338520000.0ns 0V 339320000.0ns 0V 339360000.0ns 1.95V 339760000.0ns 1.95V 339800000.0ns 0V 340600000.0ns 0V 340640000.0ns 0V 341040000.0ns 0V 341080000.0ns 0V 341880000.0ns 0V 341920000.0ns 0V 342320000.0ns 0V 342360000.0ns 0V 343160000.0ns 0V 343200000.0ns 1.95V 343600000.0ns 1.95V 343640000.0ns 0V 344440000.0ns 0V 344480000.0ns 0V 344880000.0ns 0V 344920000.0ns 0V 345720000.0ns 0V 345760000.0ns 0V 346160000.0ns 0V 346200000.0ns 0V 347000000.0ns 0V 347040000.0ns 1.95V 347440000.0ns 1.95V 347480000.0ns 0V 348280000.0ns 0V 348320000.0ns 0V 348720000.0ns 0V 348760000.0ns 0V 349560000.0ns 0V 349600000.0ns 0V 350000000.0ns 0V 350040000.0ns 0V 350840000.0ns 0V 350880000.0ns 1.95V 351280000.0ns 1.95V 351320000.0ns 0V 352120000.0ns 0V 352160000.0ns 0V 352560000.0ns 0V 352600000.0ns 0V 353400000.0ns 0V 353440000.0ns 0V 353840000.0ns 0V 353880000.0ns 0V 354680000.0ns 0V 354720000.0ns 1.95V 355120000.0ns 1.95V 355160000.0ns 0V 355960000.0ns 0V 356000000.0ns 0V 356400000.0ns 0V 356440000.0ns 0V 357240000.0ns 0V 357280000.0ns 0V 357680000.0ns 0V 357720000.0ns 0V 358520000.0ns 0V 358560000.0ns 1.95V 358960000.0ns 1.95V 359000000.0ns 0V 359800000.0ns 0V 359840000.0ns 0V 360240000.0ns 0V 360280000.0ns 0V 361080000.0ns 0V 361120000.0ns 0V 361520000.0ns 0V 361560000.0ns 0V 362360000.0ns 0V 362400000.0ns 1.95V 362800000.0ns 1.95V 362840000.0ns 0V 363640000.0ns 0V 363680000.0ns 0V 364080000.0ns 0V 364120000.0ns 0V 364920000.0ns 0V 364960000.0ns 0V 365360000.0ns 0V 365400000.0ns 0V 366200000.0ns 0V 366240000.0ns 1.95V 366640000.0ns 1.95V 366680000.0ns 0V 367480000.0ns 0V 367520000.0ns 0V 367920000.0ns 0V 367960000.0ns 0V 368760000.0ns 0V 368800000.0ns 0V 369200000.0ns 0V 369240000.0ns 0V 370040000.0ns 0V 370080000.0ns 1.95V 370480000.0ns 1.95V 370520000.0ns 0V 371320000.0ns 0V 371360000.0ns 0V 371760000.0ns 0V 371800000.0ns 0V 372600000.0ns 0V 372640000.0ns 0V 373040000.0ns 0V 373080000.0ns 0V 373880000.0ns 0V 373920000.0ns 1.95V 374320000.0ns 1.95V 374360000.0ns 0V 375160000.0ns 0V 375200000.0ns 0V 375600000.0ns 0V 375640000.0ns 0V 376440000.0ns 0V 376480000.0ns 0V 376880000.0ns 0V 376920000.0ns 0V 377720000.0ns 0V 377760000.0ns 1.95V 378160000.0ns 1.95V 378200000.0ns 0V 379000000.0ns 0V 379040000.0ns 0V 379440000.0ns 0V 379480000.0ns 0V 380280000.0ns 0V 380320000.0ns 0V 380720000.0ns 0V 380760000.0ns 0V 381560000.0ns 0V 381600000.0ns 1.95V 382000000.0ns 1.95V 382040000.0ns 0V 382840000.0ns 0V 382880000.0ns 0V 383280000.0ns 0V 383320000.0ns 0V 384120000.0ns 0V 384160000.0ns 0V 384560000.0ns 0V 384600000.0ns 0V 385400000.0ns 0V 385440000.0ns 1.95V 385840000.0ns 1.95V 385880000.0ns 0V 386680000.0ns 0V 386720000.0ns 0V 387120000.0ns 0V 387160000.0ns 0V 387960000.0ns 0V 388000000.0ns 0V 388400000.0ns 0V 388440000.0ns 0V 389240000.0ns 0V 389280000.0ns 1.95V 389680000.0ns 1.95V 389720000.0ns 0V 390520000.0ns 0V 390560000.0ns 0V 390960000.0ns 0V 391000000.0ns 0V)
VNUDGED_OUTER NUDGED_OUTER 0 PWL(0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0V 8400000.0ns 0V 8440000.0ns 0V 8920000.0ns 0V 8960000.0ns 1.95V 9680000.0ns 1.95V 9720000.0ns 0V 10200000.0ns 0V 10240000.0ns 0V 10960000.0ns 0V 11000000.0ns 0V 11480000.0ns 0V 11520000.0ns 0V 12240000.0ns 0V 12280000.0ns 0V 12760000.0ns 0V 12800000.0ns 1.95V 13520000.0ns 1.95V 13560000.0ns 0V 14040000.0ns 0V 14080000.0ns 0V 14800000.0ns 0V 14840000.0ns 0V 15320000.0ns 0V 15360000.0ns 0V 16080000.0ns 0V 16120000.0ns 0V 16600000.0ns 0V 16640000.0ns 1.95V 17360000.0ns 1.95V 17400000.0ns 0V 17880000.0ns 0V 17920000.0ns 0V 18640000.0ns 0V 18680000.0ns 0V 19160000.0ns 0V 19200000.0ns 0V 19920000.0ns 0V 19960000.0ns 0V 20440000.0ns 0V 20480000.0ns 1.95V 21200000.0ns 1.95V 21240000.0ns 0V 21720000.0ns 0V 21760000.0ns 0V 22480000.0ns 0V 22520000.0ns 0V 23000000.0ns 0V 23040000.0ns 0V 23760000.0ns 0V 23800000.0ns 0V 24280000.0ns 0V 24320000.0ns 1.95V 25040000.0ns 1.95V 25080000.0ns 0V 25560000.0ns 0V 25600000.0ns 0V 26320000.0ns 0V 26360000.0ns 0V 26840000.0ns 0V 26880000.0ns 0V 27600000.0ns 0V 27640000.0ns 0V 28120000.0ns 0V 28160000.0ns 1.95V 28880000.0ns 1.95V 28920000.0ns 0V 29400000.0ns 0V 29440000.0ns 0V 30160000.0ns 0V 30200000.0ns 0V 30680000.0ns 0V 30720000.0ns 0V 31440000.0ns 0V 31480000.0ns 0V 31960000.0ns 0V 32000000.0ns 1.95V 32720000.0ns 1.95V 32760000.0ns 0V 33240000.0ns 0V 33280000.0ns 0V 34000000.0ns 0V 34040000.0ns 0V 34520000.0ns 0V 34560000.0ns 0V 35280000.0ns 0V 35320000.0ns 0V 35800000.0ns 0V 35840000.0ns 1.95V 36560000.0ns 1.95V 36600000.0ns 0V 37080000.0ns 0V 37120000.0ns 0V 37840000.0ns 0V 37880000.0ns 0V 38360000.0ns 0V 38400000.0ns 0V 39120000.0ns 0V 39160000.0ns 0V 39640000.0ns 0V 39680000.0ns 1.95V 40400000.0ns 1.95V 40440000.0ns 0V 40920000.0ns 0V 40960000.0ns 0V 41680000.0ns 0V 41720000.0ns 0V 42200000.0ns 0V 42240000.0ns 0V 42960000.0ns 0V 43000000.0ns 0V 43480000.0ns 0V 43520000.0ns 1.95V 44240000.0ns 1.95V 44280000.0ns 0V 44760000.0ns 0V 44800000.0ns 0V 45520000.0ns 0V 45560000.0ns 0V 46040000.0ns 0V 46080000.0ns 0V 46800000.0ns 0V 46840000.0ns 0V 47320000.0ns 0V 47360000.0ns 1.95V 48080000.0ns 1.95V 48120000.0ns 0V 48600000.0ns 0V 48640000.0ns 0V 49360000.0ns 0V 49400000.0ns 0V 49880000.0ns 0V 49920000.0ns 0V 50640000.0ns 0V 50680000.0ns 0V 51160000.0ns 0V 51200000.0ns 1.95V 51920000.0ns 1.95V 51960000.0ns 0V 52440000.0ns 0V 52480000.0ns 0V 53200000.0ns 0V 53240000.0ns 0V 53720000.0ns 0V 53760000.0ns 0V 54480000.0ns 0V 54520000.0ns 0V 55000000.0ns 0V 55040000.0ns 1.95V 55760000.0ns 1.95V 55800000.0ns 0V 56280000.0ns 0V 56320000.0ns 0V 57040000.0ns 0V 57080000.0ns 0V 57560000.0ns 0V 57600000.0ns 0V 58320000.0ns 0V 58360000.0ns 0V 58840000.0ns 0V 58880000.0ns 1.95V 59600000.0ns 1.95V 59640000.0ns 0V 60120000.0ns 0V 60160000.0ns 0V 60880000.0ns 0V 60920000.0ns 0V 61400000.0ns 0V 61440000.0ns 0V 62160000.0ns 0V 62200000.0ns 0V 62680000.0ns 0V 62720000.0ns 1.95V 63440000.0ns 1.95V 63480000.0ns 0V 63960000.0ns 0V 64000000.0ns 0V 64720000.0ns 0V 64760000.0ns 0V 65240000.0ns 0V 65280000.0ns 0V 66000000.0ns 0V 66040000.0ns 0V 66520000.0ns 0V 66560000.0ns 1.95V 67280000.0ns 1.95V 67320000.0ns 0V 67800000.0ns 0V 67840000.0ns 0V 68560000.0ns 0V 68600000.0ns 0V 69080000.0ns 0V 69120000.0ns 0V 69840000.0ns 0V 69880000.0ns 0V 70360000.0ns 0V 70400000.0ns 1.95V 71120000.0ns 1.95V 71160000.0ns 0V 71640000.0ns 0V 71680000.0ns 0V 72400000.0ns 0V 72440000.0ns 0V 72920000.0ns 0V 72960000.0ns 0V 73680000.0ns 0V 73720000.0ns 0V 74200000.0ns 0V 74240000.0ns 1.95V 74960000.0ns 1.95V 75000000.0ns 0V 75480000.0ns 0V 75520000.0ns 0V 76240000.0ns 0V 76280000.0ns 0V 76760000.0ns 0V 76800000.0ns 0V 77520000.0ns 0V 77560000.0ns 0V 78040000.0ns 0V 78080000.0ns 1.95V 78800000.0ns 1.95V 78840000.0ns 0V 79320000.0ns 0V 79360000.0ns 0V 80080000.0ns 0V 80120000.0ns 0V 80600000.0ns 0V 80640000.0ns 0V 81360000.0ns 0V 81400000.0ns 0V 81880000.0ns 0V 81920000.0ns 1.95V 82640000.0ns 1.95V 82680000.0ns 0V 83160000.0ns 0V 83200000.0ns 0V 83920000.0ns 0V 83960000.0ns 0V 84440000.0ns 0V 84480000.0ns 0V 85200000.0ns 0V 85240000.0ns 0V 85720000.0ns 0V 85760000.0ns 1.95V 86480000.0ns 1.95V 86520000.0ns 0V 87000000.0ns 0V 87040000.0ns 0V 87760000.0ns 0V 87800000.0ns 0V 88280000.0ns 0V 88320000.0ns 0V 89040000.0ns 0V 89080000.0ns 0V 89560000.0ns 0V 89600000.0ns 1.95V 90320000.0ns 1.95V 90360000.0ns 0V 90840000.0ns 0V 90880000.0ns 0V 91600000.0ns 0V 91640000.0ns 0V 92120000.0ns 0V 92160000.0ns 0V 92880000.0ns 0V 92920000.0ns 0V 93400000.0ns 0V 93440000.0ns 1.95V 94160000.0ns 1.95V 94200000.0ns 0V 94680000.0ns 0V 94720000.0ns 0V 95440000.0ns 0V 95480000.0ns 0V 95960000.0ns 0V 96000000.0ns 0V 96720000.0ns 0V 96760000.0ns 0V 97240000.0ns 0V 97280000.0ns 1.95V 98000000.0ns 1.95V 98040000.0ns 0V 98520000.0ns 0V 98560000.0ns 0V 99280000.0ns 0V 99320000.0ns 0V 99800000.0ns 0V 99840000.0ns 0V 100560000.0ns 0V 100600000.0ns 0V 101080000.0ns 0V 101120000.0ns 1.95V 101840000.0ns 1.95V 101880000.0ns 0V 102360000.0ns 0V 102400000.0ns 0V 103120000.0ns 0V 103160000.0ns 0V 103640000.0ns 0V 103680000.0ns 0V 104400000.0ns 0V 104440000.0ns 0V 104920000.0ns 0V 104960000.0ns 1.95V 105680000.0ns 1.95V 105720000.0ns 0V 106200000.0ns 0V 106240000.0ns 0V 106960000.0ns 0V 107000000.0ns 0V 107480000.0ns 0V 107520000.0ns 0V 108240000.0ns 0V 108280000.0ns 0V 108760000.0ns 0V 108800000.0ns 1.95V 109520000.0ns 1.95V 109560000.0ns 0V 110040000.0ns 0V 110080000.0ns 0V 110800000.0ns 0V 110840000.0ns 0V 111320000.0ns 0V 111360000.0ns 0V 112080000.0ns 0V 112120000.0ns 0V 112600000.0ns 0V 112640000.0ns 1.95V 113360000.0ns 1.95V 113400000.0ns 0V 113880000.0ns 0V 113920000.0ns 0V 114640000.0ns 0V 114680000.0ns 0V 115160000.0ns 0V 115200000.0ns 0V 115920000.0ns 0V 115960000.0ns 0V 116440000.0ns 0V 116480000.0ns 1.95V 117200000.0ns 1.95V 117240000.0ns 0V 117720000.0ns 0V 117760000.0ns 0V 118480000.0ns 0V 118520000.0ns 0V 119000000.0ns 0V 119040000.0ns 0V 119760000.0ns 0V 119800000.0ns 0V 120280000.0ns 0V 120320000.0ns 1.95V 121040000.0ns 1.95V 121080000.0ns 0V 121560000.0ns 0V 121600000.0ns 0V 122320000.0ns 0V 122360000.0ns 0V 122840000.0ns 0V 122880000.0ns 0V 123600000.0ns 0V 123640000.0ns 0V 124120000.0ns 0V 124160000.0ns 1.95V 124880000.0ns 1.95V 124920000.0ns 0V 125400000.0ns 0V 125440000.0ns 0V 126160000.0ns 0V 126200000.0ns 0V 126680000.0ns 0V 126720000.0ns 0V 127440000.0ns 0V 127480000.0ns 0V 127960000.0ns 0V 128000000.0ns 1.95V 128720000.0ns 1.95V 128760000.0ns 0V 129240000.0ns 0V 129280000.0ns 0V 130000000.0ns 0V 130040000.0ns 0V 130520000.0ns 0V 130560000.0ns 0V 131280000.0ns 0V 131320000.0ns 0V 131800000.0ns 0V 131840000.0ns 1.95V 132560000.0ns 1.95V 132600000.0ns 0V 133080000.0ns 0V 133120000.0ns 0V 133840000.0ns 0V 133880000.0ns 0V 134360000.0ns 0V 134400000.0ns 0V 135120000.0ns 0V 135160000.0ns 0V 135640000.0ns 0V 135680000.0ns 1.95V 136400000.0ns 1.95V 136440000.0ns 0V 136920000.0ns 0V 136960000.0ns 0V 137680000.0ns 0V 137720000.0ns 0V 138200000.0ns 0V 138240000.0ns 0V 138960000.0ns 0V 139000000.0ns 0V 139480000.0ns 0V 139520000.0ns 1.95V 140240000.0ns 1.95V 140280000.0ns 0V 140760000.0ns 0V 140800000.0ns 0V 141520000.0ns 0V 141560000.0ns 0V 142040000.0ns 0V 142080000.0ns 0V 142800000.0ns 0V 142840000.0ns 0V 143320000.0ns 0V 143360000.0ns 1.95V 144080000.0ns 1.95V 144120000.0ns 0V 144600000.0ns 0V 144640000.0ns 0V 145360000.0ns 0V 145400000.0ns 0V 145880000.0ns 0V 145920000.0ns 0V 146640000.0ns 0V 146680000.0ns 0V 147160000.0ns 0V 147200000.0ns 1.95V 147920000.0ns 1.95V 147960000.0ns 0V 148440000.0ns 0V 148480000.0ns 0V 149200000.0ns 0V 149240000.0ns 0V 149720000.0ns 0V 149760000.0ns 0V 150480000.0ns 0V 150520000.0ns 0V 151000000.0ns 0V 151040000.0ns 1.95V 151760000.0ns 1.95V 151800000.0ns 0V 152280000.0ns 0V 152320000.0ns 0V 153040000.0ns 0V 153080000.0ns 0V 153560000.0ns 0V 153600000.0ns 0V 154320000.0ns 0V 154360000.0ns 0V 154840000.0ns 0V 154880000.0ns 1.95V 155600000.0ns 1.95V 155640000.0ns 0V 156120000.0ns 0V 156160000.0ns 0V 156880000.0ns 0V 156920000.0ns 0V 157400000.0ns 0V 157440000.0ns 0V 158160000.0ns 0V 158200000.0ns 0V 158680000.0ns 0V 158720000.0ns 1.95V 159440000.0ns 1.95V 159480000.0ns 0V 159960000.0ns 0V 160000000.0ns 0V 160720000.0ns 0V 160760000.0ns 0V 161240000.0ns 0V 161280000.0ns 0V 162000000.0ns 0V 162040000.0ns 0V 162520000.0ns 0V 162560000.0ns 1.95V 163280000.0ns 1.95V 163320000.0ns 0V 163800000.0ns 0V 163840000.0ns 0V 164560000.0ns 0V 164600000.0ns 0V 165080000.0ns 0V 165120000.0ns 0V 165840000.0ns 0V 165880000.0ns 0V 166360000.0ns 0V 166400000.0ns 1.95V 167120000.0ns 1.95V 167160000.0ns 0V 167640000.0ns 0V 167680000.0ns 0V 168400000.0ns 0V 168440000.0ns 0V 168920000.0ns 0V 168960000.0ns 0V 169680000.0ns 0V 169720000.0ns 0V 170200000.0ns 0V 170240000.0ns 1.95V 170960000.0ns 1.95V 171000000.0ns 0V 171480000.0ns 0V 171520000.0ns 0V 172240000.0ns 0V 172280000.0ns 0V 172760000.0ns 0V 172800000.0ns 0V 173520000.0ns 0V 173560000.0ns 0V 174040000.0ns 0V 174080000.0ns 1.95V 174800000.0ns 1.95V 174840000.0ns 0V 175320000.0ns 0V 175360000.0ns 0V 176080000.0ns 0V 176120000.0ns 0V 176600000.0ns 0V 176640000.0ns 0V 177360000.0ns 0V 177400000.0ns 0V 177880000.0ns 0V 177920000.0ns 1.95V 178640000.0ns 1.95V 178680000.0ns 0V 179160000.0ns 0V 179200000.0ns 0V 179920000.0ns 0V 179960000.0ns 0V 180440000.0ns 0V 180480000.0ns 0V 181200000.0ns 0V 181240000.0ns 0V 181720000.0ns 0V 181760000.0ns 1.95V 182480000.0ns 1.95V 182520000.0ns 0V 183000000.0ns 0V 183040000.0ns 0V 183760000.0ns 0V 183800000.0ns 0V 184280000.0ns 0V 184320000.0ns 0V 185040000.0ns 0V 185080000.0ns 0V 185560000.0ns 0V 185600000.0ns 1.95V 186320000.0ns 1.95V 186360000.0ns 0V 186840000.0ns 0V 186880000.0ns 0V 187600000.0ns 0V 187640000.0ns 0V 188120000.0ns 0V 188160000.0ns 0V 188880000.0ns 0V 188920000.0ns 0V 189400000.0ns 0V 189440000.0ns 1.95V 190160000.0ns 1.95V 190200000.0ns 0V 190680000.0ns 0V 190720000.0ns 0V 191440000.0ns 0V 191480000.0ns 0V 191960000.0ns 0V 192000000.0ns 0V 192720000.0ns 0V 192760000.0ns 0V 193240000.0ns 0V 193280000.0ns 1.95V 194000000.0ns 1.95V 194040000.0ns 0V 194520000.0ns 0V 194560000.0ns 0V 195280000.0ns 0V 195320000.0ns 0V 195800000.0ns 0V 195840000.0ns 0V 196560000.0ns 0V 196600000.0ns 0V 197080000.0ns 0V 197120000.0ns 1.95V 197840000.0ns 1.95V 197880000.0ns 0V 198360000.0ns 0V 198400000.0ns 0V 199120000.0ns 0V 199160000.0ns 0V 199640000.0ns 0V 199680000.0ns 0V 200400000.0ns 0V 200440000.0ns 0V 200920000.0ns 0V 200960000.0ns 1.95V 201680000.0ns 1.95V 201720000.0ns 0V 202200000.0ns 0V 202240000.0ns 0V 202960000.0ns 0V 203000000.0ns 0V 203480000.0ns 0V 203520000.0ns 0V 204240000.0ns 0V 204280000.0ns 0V 204760000.0ns 0V 204800000.0ns 1.95V 205520000.0ns 1.95V 205560000.0ns 0V 206040000.0ns 0V 206080000.0ns 0V 206800000.0ns 0V 206840000.0ns 0V 207320000.0ns 0V 207360000.0ns 0V 208080000.0ns 0V 208120000.0ns 0V 208600000.0ns 0V 208640000.0ns 1.95V 209360000.0ns 1.95V 209400000.0ns 0V 209880000.0ns 0V 209920000.0ns 0V 210640000.0ns 0V 210680000.0ns 0V 211160000.0ns 0V 211200000.0ns 0V 211920000.0ns 0V 211960000.0ns 0V 212440000.0ns 0V 212480000.0ns 1.95V 213200000.0ns 1.95V 213240000.0ns 0V 213720000.0ns 0V 213760000.0ns 0V 214480000.0ns 0V 214520000.0ns 0V 215000000.0ns 0V 215040000.0ns 0V 215760000.0ns 0V 215800000.0ns 0V 216280000.0ns 0V 216320000.0ns 1.95V 217040000.0ns 1.95V 217080000.0ns 0V 217560000.0ns 0V 217600000.0ns 0V 218320000.0ns 0V 218360000.0ns 0V 218840000.0ns 0V 218880000.0ns 0V 219600000.0ns 0V 219640000.0ns 0V 220120000.0ns 0V 220160000.0ns 1.95V 220880000.0ns 1.95V 220920000.0ns 0V 221400000.0ns 0V 221440000.0ns 0V 222160000.0ns 0V 222200000.0ns 0V 222680000.0ns 0V 222720000.0ns 0V 223440000.0ns 0V 223480000.0ns 0V 223960000.0ns 0V 224000000.0ns 1.95V 224720000.0ns 1.95V 224760000.0ns 0V 225240000.0ns 0V 225280000.0ns 0V 226000000.0ns 0V 226040000.0ns 0V 226520000.0ns 0V 226560000.0ns 0V 227280000.0ns 0V 227320000.0ns 0V 227800000.0ns 0V 227840000.0ns 1.95V 228560000.0ns 1.95V 228600000.0ns 0V 229080000.0ns 0V 229120000.0ns 0V 229840000.0ns 0V 229880000.0ns 0V 230360000.0ns 0V 230400000.0ns 0V 231120000.0ns 0V 231160000.0ns 0V 231640000.0ns 0V 231680000.0ns 1.95V 232400000.0ns 1.95V 232440000.0ns 0V 232920000.0ns 0V 232960000.0ns 0V 233680000.0ns 0V 233720000.0ns 0V 234200000.0ns 0V 234240000.0ns 0V 234960000.0ns 0V 235000000.0ns 0V 235480000.0ns 0V 235520000.0ns 1.95V 236240000.0ns 1.95V 236280000.0ns 0V 236760000.0ns 0V 236800000.0ns 0V 237520000.0ns 0V 237560000.0ns 0V 238040000.0ns 0V 238080000.0ns 0V 238800000.0ns 0V 238840000.0ns 0V 239320000.0ns 0V 239360000.0ns 1.95V 240080000.0ns 1.95V 240120000.0ns 0V 240600000.0ns 0V 240640000.0ns 0V 241360000.0ns 0V 241400000.0ns 0V 241880000.0ns 0V 241920000.0ns 0V 242640000.0ns 0V 242680000.0ns 0V 243160000.0ns 0V 243200000.0ns 1.95V 243920000.0ns 1.95V 243960000.0ns 0V 244440000.0ns 0V 244480000.0ns 0V 245200000.0ns 0V 245240000.0ns 0V 245720000.0ns 0V 245760000.0ns 0V 246480000.0ns 0V 246520000.0ns 0V 247000000.0ns 0V 247040000.0ns 1.95V 247760000.0ns 1.95V 247800000.0ns 0V 248280000.0ns 0V 248320000.0ns 0V 249040000.0ns 0V 249080000.0ns 0V 249560000.0ns 0V 249600000.0ns 0V 250320000.0ns 0V 250360000.0ns 0V 250840000.0ns 0V 250880000.0ns 1.95V 251600000.0ns 1.95V 251640000.0ns 0V 252120000.0ns 0V 252160000.0ns 0V 252880000.0ns 0V 252920000.0ns 0V 253400000.0ns 0V 253440000.0ns 0V 254160000.0ns 0V 254200000.0ns 0V 254680000.0ns 0V 254720000.0ns 1.95V 255440000.0ns 1.95V 255480000.0ns 0V 255960000.0ns 0V 256000000.0ns 0V 256720000.0ns 0V 256760000.0ns 0V 257240000.0ns 0V 257280000.0ns 0V 258000000.0ns 0V 258040000.0ns 0V 258520000.0ns 0V 258560000.0ns 1.95V 259280000.0ns 1.95V 259320000.0ns 0V 259800000.0ns 0V 259840000.0ns 0V 260560000.0ns 0V 260600000.0ns 0V 261080000.0ns 0V 261120000.0ns 0V 261840000.0ns 0V 261880000.0ns 0V 262360000.0ns 0V 262400000.0ns 1.95V 263120000.0ns 1.95V 263160000.0ns 0V 263640000.0ns 0V 263680000.0ns 0V 264400000.0ns 0V 264440000.0ns 0V 264920000.0ns 0V 264960000.0ns 0V 265680000.0ns 0V 265720000.0ns 0V 266200000.0ns 0V 266240000.0ns 1.95V 266960000.0ns 1.95V 267000000.0ns 0V 267480000.0ns 0V 267520000.0ns 0V 268240000.0ns 0V 268280000.0ns 0V 268760000.0ns 0V 268800000.0ns 0V 269520000.0ns 0V 269560000.0ns 0V 270040000.0ns 0V 270080000.0ns 1.95V 270800000.0ns 1.95V 270840000.0ns 0V 271320000.0ns 0V 271360000.0ns 0V 272080000.0ns 0V 272120000.0ns 0V 272600000.0ns 0V 272640000.0ns 0V 273360000.0ns 0V 273400000.0ns 0V 273880000.0ns 0V 273920000.0ns 1.95V 274640000.0ns 1.95V 274680000.0ns 0V 275160000.0ns 0V 275200000.0ns 0V 275920000.0ns 0V 275960000.0ns 0V 276440000.0ns 0V 276480000.0ns 0V 277200000.0ns 0V 277240000.0ns 0V 277720000.0ns 0V 277760000.0ns 1.95V 278480000.0ns 1.95V 278520000.0ns 0V 279000000.0ns 0V 279040000.0ns 0V 279760000.0ns 0V 279800000.0ns 0V 280280000.0ns 0V 280320000.0ns 0V 281040000.0ns 0V 281080000.0ns 0V 281560000.0ns 0V 281600000.0ns 1.95V 282320000.0ns 1.95V 282360000.0ns 0V 282840000.0ns 0V 282880000.0ns 0V 283600000.0ns 0V 283640000.0ns 0V 284120000.0ns 0V 284160000.0ns 0V 284880000.0ns 0V 284920000.0ns 0V 285400000.0ns 0V 285440000.0ns 1.95V 286160000.0ns 1.95V 286200000.0ns 0V 286680000.0ns 0V 286720000.0ns 0V 287440000.0ns 0V 287480000.0ns 0V 287960000.0ns 0V 288000000.0ns 0V 288720000.0ns 0V 288760000.0ns 0V 289240000.0ns 0V 289280000.0ns 1.95V 290000000.0ns 1.95V 290040000.0ns 0V 290520000.0ns 0V 290560000.0ns 0V 291280000.0ns 0V 291320000.0ns 0V 291800000.0ns 0V 291840000.0ns 0V 292560000.0ns 0V 292600000.0ns 0V 293080000.0ns 0V 293120000.0ns 1.95V 293840000.0ns 1.95V 293880000.0ns 0V 294360000.0ns 0V 294400000.0ns 0V 295120000.0ns 0V 295160000.0ns 0V 295640000.0ns 0V 295680000.0ns 0V 296400000.0ns 0V 296440000.0ns 0V 296920000.0ns 0V 296960000.0ns 1.95V 297680000.0ns 1.95V 297720000.0ns 0V 298200000.0ns 0V 298240000.0ns 0V 298960000.0ns 0V 299000000.0ns 0V 299480000.0ns 0V 299520000.0ns 0V 300240000.0ns 0V 300280000.0ns 0V 300760000.0ns 0V 300800000.0ns 1.95V 301520000.0ns 1.95V 301560000.0ns 0V 302040000.0ns 0V 302080000.0ns 0V 302800000.0ns 0V 302840000.0ns 0V 303320000.0ns 0V 303360000.0ns 0V 304080000.0ns 0V 304120000.0ns 0V 304600000.0ns 0V 304640000.0ns 1.95V 305360000.0ns 1.95V 305400000.0ns 0V 305880000.0ns 0V 305920000.0ns 0V 306640000.0ns 0V 306680000.0ns 0V 307160000.0ns 0V 307200000.0ns 0V 307920000.0ns 0V 307960000.0ns 0V 308440000.0ns 0V 308480000.0ns 1.95V 309200000.0ns 1.95V 309240000.0ns 0V 309720000.0ns 0V 309760000.0ns 0V 310480000.0ns 0V 310520000.0ns 0V 311000000.0ns 0V 311040000.0ns 0V 311760000.0ns 0V 311800000.0ns 0V 312280000.0ns 0V 312320000.0ns 1.95V 313040000.0ns 1.95V 313080000.0ns 0V 313560000.0ns 0V 313600000.0ns 0V 314320000.0ns 0V 314360000.0ns 0V 314840000.0ns 0V 314880000.0ns 0V 315600000.0ns 0V 315640000.0ns 0V 316120000.0ns 0V 316160000.0ns 1.95V 316880000.0ns 1.95V 316920000.0ns 0V 317400000.0ns 0V 317440000.0ns 0V 318160000.0ns 0V 318200000.0ns 0V 318680000.0ns 0V 318720000.0ns 0V 319440000.0ns 0V 319480000.0ns 0V 319960000.0ns 0V 320000000.0ns 1.95V 320720000.0ns 1.95V 320760000.0ns 0V 321240000.0ns 0V 321280000.0ns 0V 322000000.0ns 0V 322040000.0ns 0V 322520000.0ns 0V 322560000.0ns 0V 323280000.0ns 0V 323320000.0ns 0V 323800000.0ns 0V 323840000.0ns 1.95V 324560000.0ns 1.95V 324600000.0ns 0V 325080000.0ns 0V 325120000.0ns 0V 325840000.0ns 0V 325880000.0ns 0V 326360000.0ns 0V 326400000.0ns 0V 327120000.0ns 0V 327160000.0ns 0V 327640000.0ns 0V 327680000.0ns 1.95V 328400000.0ns 1.95V 328440000.0ns 0V 328920000.0ns 0V 328960000.0ns 0V 329680000.0ns 0V 329720000.0ns 0V 330200000.0ns 0V 330240000.0ns 0V 330960000.0ns 0V 331000000.0ns 0V 331480000.0ns 0V 331520000.0ns 1.95V 332240000.0ns 1.95V 332280000.0ns 0V 332760000.0ns 0V 332800000.0ns 0V 333520000.0ns 0V 333560000.0ns 0V 334040000.0ns 0V 334080000.0ns 0V 334800000.0ns 0V 334840000.0ns 0V 335320000.0ns 0V 335360000.0ns 1.95V 336080000.0ns 1.95V 336120000.0ns 0V 336600000.0ns 0V 336640000.0ns 0V 337360000.0ns 0V 337400000.0ns 0V 337880000.0ns 0V 337920000.0ns 0V 338640000.0ns 0V 338680000.0ns 0V 339160000.0ns 0V 339200000.0ns 1.95V 339920000.0ns 1.95V 339960000.0ns 0V 340440000.0ns 0V 340480000.0ns 0V 341200000.0ns 0V 341240000.0ns 0V 341720000.0ns 0V 341760000.0ns 0V 342480000.0ns 0V 342520000.0ns 0V 343000000.0ns 0V 343040000.0ns 1.95V 343760000.0ns 1.95V 343800000.0ns 0V 344280000.0ns 0V 344320000.0ns 0V 345040000.0ns 0V 345080000.0ns 0V 345560000.0ns 0V 345600000.0ns 0V 346320000.0ns 0V 346360000.0ns 0V 346840000.0ns 0V 346880000.0ns 1.95V 347600000.0ns 1.95V 347640000.0ns 0V 348120000.0ns 0V 348160000.0ns 0V 348880000.0ns 0V 348920000.0ns 0V 349400000.0ns 0V 349440000.0ns 0V 350160000.0ns 0V 350200000.0ns 0V 350680000.0ns 0V 350720000.0ns 1.95V 351440000.0ns 1.95V 351480000.0ns 0V 351960000.0ns 0V 352000000.0ns 0V 352720000.0ns 0V 352760000.0ns 0V 353240000.0ns 0V 353280000.0ns 0V 354000000.0ns 0V 354040000.0ns 0V 354520000.0ns 0V 354560000.0ns 1.95V 355280000.0ns 1.95V 355320000.0ns 0V 355800000.0ns 0V 355840000.0ns 0V 356560000.0ns 0V 356600000.0ns 0V 357080000.0ns 0V 357120000.0ns 0V 357840000.0ns 0V 357880000.0ns 0V 358360000.0ns 0V 358400000.0ns 1.95V 359120000.0ns 1.95V 359160000.0ns 0V 359640000.0ns 0V 359680000.0ns 0V 360400000.0ns 0V 360440000.0ns 0V 360920000.0ns 0V 360960000.0ns 0V 361680000.0ns 0V 361720000.0ns 0V 362200000.0ns 0V 362240000.0ns 1.95V 362960000.0ns 1.95V 363000000.0ns 0V 363480000.0ns 0V 363520000.0ns 0V 364240000.0ns 0V 364280000.0ns 0V 364760000.0ns 0V 364800000.0ns 0V 365520000.0ns 0V 365560000.0ns 0V 366040000.0ns 0V 366080000.0ns 1.95V 366800000.0ns 1.95V 366840000.0ns 0V 367320000.0ns 0V 367360000.0ns 0V 368080000.0ns 0V 368120000.0ns 0V 368600000.0ns 0V 368640000.0ns 0V 369360000.0ns 0V 369400000.0ns 0V 369880000.0ns 0V 369920000.0ns 1.95V 370640000.0ns 1.95V 370680000.0ns 0V 371160000.0ns 0V 371200000.0ns 0V 371920000.0ns 0V 371960000.0ns 0V 372440000.0ns 0V 372480000.0ns 0V 373200000.0ns 0V 373240000.0ns 0V 373720000.0ns 0V 373760000.0ns 1.95V 374480000.0ns 1.95V 374520000.0ns 0V 375000000.0ns 0V 375040000.0ns 0V 375760000.0ns 0V 375800000.0ns 0V 376280000.0ns 0V 376320000.0ns 0V 377040000.0ns 0V 377080000.0ns 0V 377560000.0ns 0V 377600000.0ns 1.95V 378320000.0ns 1.95V 378360000.0ns 0V 378840000.0ns 0V 378880000.0ns 0V 379600000.0ns 0V 379640000.0ns 0V 380120000.0ns 0V 380160000.0ns 0V 380880000.0ns 0V 380920000.0ns 0V 381400000.0ns 0V 381440000.0ns 1.95V 382160000.0ns 1.95V 382200000.0ns 0V 382680000.0ns 0V 382720000.0ns 0V 383440000.0ns 0V 383480000.0ns 0V 383960000.0ns 0V 384000000.0ns 0V 384720000.0ns 0V 384760000.0ns 0V 385240000.0ns 0V 385280000.0ns 1.95V 386000000.0ns 1.95V 386040000.0ns 0V 386520000.0ns 0V 386560000.0ns 0V 387280000.0ns 0V 387320000.0ns 0V 387800000.0ns 0V 387840000.0ns 0V 388560000.0ns 0V 388600000.0ns 0V 389080000.0ns 0V 389120000.0ns 1.95V 389840000.0ns 1.95V 389880000.0ns 0V 390360000.0ns 0V 390400000.0ns 0V 391120000.0ns 0V 391160000.0ns 0V)
VFREE FREE 0 PWL(0ns 0V 3960000.0ns 0V 7800000.0ns 0V 7840000.0ns 1.95V 8240000.0ns 1.95V 8280000.0ns 0V 9080000.0ns 0V 9120000.0ns 0V 9520000.0ns 0V 9560000.0ns 0V 10360000.0ns 0V 10400000.0ns 0V 10800000.0ns 0V 10840000.0ns 0V 11640000.0ns 0V 11680000.0ns 1.95V 12080000.0ns 1.95V 12120000.0ns 0V 12920000.0ns 0V 12960000.0ns 0V 13360000.0ns 0V 13400000.0ns 0V 14200000.0ns 0V 14240000.0ns 0V 14640000.0ns 0V 14680000.0ns 0V 15480000.0ns 0V 15520000.0ns 1.95V 15920000.0ns 1.95V 15960000.0ns 0V 16760000.0ns 0V 16800000.0ns 0V 17200000.0ns 0V 17240000.0ns 0V 18040000.0ns 0V 18080000.0ns 0V 18480000.0ns 0V 18520000.0ns 0V 19320000.0ns 0V 19360000.0ns 1.95V 19760000.0ns 1.95V 19800000.0ns 0V 20600000.0ns 0V 20640000.0ns 0V 21040000.0ns 0V 21080000.0ns 0V 21880000.0ns 0V 21920000.0ns 0V 22320000.0ns 0V 22360000.0ns 0V 23160000.0ns 0V 23200000.0ns 1.95V 23600000.0ns 1.95V 23640000.0ns 0V 24440000.0ns 0V 24480000.0ns 0V 24880000.0ns 0V 24920000.0ns 0V 25720000.0ns 0V 25760000.0ns 0V 26160000.0ns 0V 26200000.0ns 0V 27000000.0ns 0V 27040000.0ns 1.95V 27440000.0ns 1.95V 27480000.0ns 0V 28280000.0ns 0V 28320000.0ns 0V 28720000.0ns 0V 28760000.0ns 0V 29560000.0ns 0V 29600000.0ns 0V 30000000.0ns 0V 30040000.0ns 0V 30840000.0ns 0V 30880000.0ns 1.95V 31280000.0ns 1.95V 31320000.0ns 0V 32120000.0ns 0V 32160000.0ns 0V 32560000.0ns 0V 32600000.0ns 0V 33400000.0ns 0V 33440000.0ns 0V 33840000.0ns 0V 33880000.0ns 0V 34680000.0ns 0V 34720000.0ns 1.95V 35120000.0ns 1.95V 35160000.0ns 0V 35960000.0ns 0V 36000000.0ns 0V 36400000.0ns 0V 36440000.0ns 0V 37240000.0ns 0V 37280000.0ns 0V 37680000.0ns 0V 37720000.0ns 0V 38520000.0ns 0V 38560000.0ns 1.95V 38960000.0ns 1.95V 39000000.0ns 0V 39800000.0ns 0V 39840000.0ns 0V 40240000.0ns 0V 40280000.0ns 0V 41080000.0ns 0V 41120000.0ns 0V 41520000.0ns 0V 41560000.0ns 0V 42360000.0ns 0V 42400000.0ns 1.95V 42800000.0ns 1.95V 42840000.0ns 0V 43640000.0ns 0V 43680000.0ns 0V 44080000.0ns 0V 44120000.0ns 0V 44920000.0ns 0V 44960000.0ns 0V 45360000.0ns 0V 45400000.0ns 0V 46200000.0ns 0V 46240000.0ns 1.95V 46640000.0ns 1.95V 46680000.0ns 0V 47480000.0ns 0V 47520000.0ns 0V 47920000.0ns 0V 47960000.0ns 0V 48760000.0ns 0V 48800000.0ns 0V 49200000.0ns 0V 49240000.0ns 0V 50040000.0ns 0V 50080000.0ns 1.95V 50480000.0ns 1.95V 50520000.0ns 0V 51320000.0ns 0V 51360000.0ns 0V 51760000.0ns 0V 51800000.0ns 0V 52600000.0ns 0V 52640000.0ns 0V 53040000.0ns 0V 53080000.0ns 0V 53880000.0ns 0V 53920000.0ns 1.95V 54320000.0ns 1.95V 54360000.0ns 0V 55160000.0ns 0V 55200000.0ns 0V 55600000.0ns 0V 55640000.0ns 0V 56440000.0ns 0V 56480000.0ns 0V 56880000.0ns 0V 56920000.0ns 0V 57720000.0ns 0V 57760000.0ns 1.95V 58160000.0ns 1.95V 58200000.0ns 0V 59000000.0ns 0V 59040000.0ns 0V 59440000.0ns 0V 59480000.0ns 0V 60280000.0ns 0V 60320000.0ns 0V 60720000.0ns 0V 60760000.0ns 0V 61560000.0ns 0V 61600000.0ns 1.95V 62000000.0ns 1.95V 62040000.0ns 0V 62840000.0ns 0V 62880000.0ns 0V 63280000.0ns 0V 63320000.0ns 0V 64120000.0ns 0V 64160000.0ns 0V 64560000.0ns 0V 64600000.0ns 0V 65400000.0ns 0V 65440000.0ns 1.95V 65840000.0ns 1.95V 65880000.0ns 0V 66680000.0ns 0V 66720000.0ns 0V 67120000.0ns 0V 67160000.0ns 0V 67960000.0ns 0V 68000000.0ns 0V 68400000.0ns 0V 68440000.0ns 0V 69240000.0ns 0V 69280000.0ns 1.95V 69680000.0ns 1.95V 69720000.0ns 0V 70520000.0ns 0V 70560000.0ns 0V 70960000.0ns 0V 71000000.0ns 0V 71800000.0ns 0V 71840000.0ns 0V 72240000.0ns 0V 72280000.0ns 0V 73080000.0ns 0V 73120000.0ns 1.95V 73520000.0ns 1.95V 73560000.0ns 0V 74360000.0ns 0V 74400000.0ns 0V 74800000.0ns 0V 74840000.0ns 0V 75640000.0ns 0V 75680000.0ns 0V 76080000.0ns 0V 76120000.0ns 0V 76920000.0ns 0V 76960000.0ns 1.95V 77360000.0ns 1.95V 77400000.0ns 0V 78200000.0ns 0V 78240000.0ns 0V 78640000.0ns 0V 78680000.0ns 0V 79480000.0ns 0V 79520000.0ns 0V 79920000.0ns 0V 79960000.0ns 0V 80760000.0ns 0V 80800000.0ns 1.95V 81200000.0ns 1.95V 81240000.0ns 0V 82040000.0ns 0V 82080000.0ns 0V 82480000.0ns 0V 82520000.0ns 0V 83320000.0ns 0V 83360000.0ns 0V 83760000.0ns 0V 83800000.0ns 0V 84600000.0ns 0V 84640000.0ns 1.95V 85040000.0ns 1.95V 85080000.0ns 0V 85880000.0ns 0V 85920000.0ns 0V 86320000.0ns 0V 86360000.0ns 0V 87160000.0ns 0V 87200000.0ns 0V 87600000.0ns 0V 87640000.0ns 0V 88440000.0ns 0V 88480000.0ns 1.95V 88880000.0ns 1.95V 88920000.0ns 0V 89720000.0ns 0V 89760000.0ns 0V 90160000.0ns 0V 90200000.0ns 0V 91000000.0ns 0V 91040000.0ns 0V 91440000.0ns 0V 91480000.0ns 0V 92280000.0ns 0V 92320000.0ns 1.95V 92720000.0ns 1.95V 92760000.0ns 0V 93560000.0ns 0V 93600000.0ns 0V 94000000.0ns 0V 94040000.0ns 0V 94840000.0ns 0V 94880000.0ns 0V 95280000.0ns 0V 95320000.0ns 0V 96120000.0ns 0V 96160000.0ns 1.95V 96560000.0ns 1.95V 96600000.0ns 0V 97400000.0ns 0V 97440000.0ns 0V 97840000.0ns 0V 97880000.0ns 0V 98680000.0ns 0V 98720000.0ns 0V 99120000.0ns 0V 99160000.0ns 0V 99960000.0ns 0V 100000000.0ns 1.95V 100400000.0ns 1.95V 100440000.0ns 0V 101240000.0ns 0V 101280000.0ns 0V 101680000.0ns 0V 101720000.0ns 0V 102520000.0ns 0V 102560000.0ns 0V 102960000.0ns 0V 103000000.0ns 0V 103800000.0ns 0V 103840000.0ns 1.95V 104240000.0ns 1.95V 104280000.0ns 0V 105080000.0ns 0V 105120000.0ns 0V 105520000.0ns 0V 105560000.0ns 0V 106360000.0ns 0V 106400000.0ns 0V 106800000.0ns 0V 106840000.0ns 0V 107640000.0ns 0V 107680000.0ns 1.95V 108080000.0ns 1.95V 108120000.0ns 0V 108920000.0ns 0V 108960000.0ns 0V 109360000.0ns 0V 109400000.0ns 0V 110200000.0ns 0V 110240000.0ns 0V 110640000.0ns 0V 110680000.0ns 0V 111480000.0ns 0V 111520000.0ns 1.95V 111920000.0ns 1.95V 111960000.0ns 0V 112760000.0ns 0V 112800000.0ns 0V 113200000.0ns 0V 113240000.0ns 0V 114040000.0ns 0V 114080000.0ns 0V 114480000.0ns 0V 114520000.0ns 0V 115320000.0ns 0V 115360000.0ns 1.95V 115760000.0ns 1.95V 115800000.0ns 0V 116600000.0ns 0V 116640000.0ns 0V 117040000.0ns 0V 117080000.0ns 0V 117880000.0ns 0V 117920000.0ns 0V 118320000.0ns 0V 118360000.0ns 0V 119160000.0ns 0V 119200000.0ns 1.95V 119600000.0ns 1.95V 119640000.0ns 0V 120440000.0ns 0V 120480000.0ns 0V 120880000.0ns 0V 120920000.0ns 0V 121720000.0ns 0V 121760000.0ns 0V 122160000.0ns 0V 122200000.0ns 0V 123000000.0ns 0V 123040000.0ns 1.95V 123440000.0ns 1.95V 123480000.0ns 0V 124280000.0ns 0V 124320000.0ns 0V 124720000.0ns 0V 124760000.0ns 0V 125560000.0ns 0V 125600000.0ns 0V 126000000.0ns 0V 126040000.0ns 0V 126840000.0ns 0V 126880000.0ns 1.95V 127280000.0ns 1.95V 127320000.0ns 0V 128120000.0ns 0V 128160000.0ns 0V 128560000.0ns 0V 128600000.0ns 0V 129400000.0ns 0V 129440000.0ns 0V 129840000.0ns 0V 129880000.0ns 0V 130680000.0ns 0V 130720000.0ns 1.95V 131120000.0ns 1.95V 131160000.0ns 0V 131960000.0ns 0V 132000000.0ns 0V 132400000.0ns 0V 132440000.0ns 0V 133240000.0ns 0V 133280000.0ns 0V 133680000.0ns 0V 133720000.0ns 0V 134520000.0ns 0V 134560000.0ns 1.95V 134960000.0ns 1.95V 135000000.0ns 0V 135800000.0ns 0V 135840000.0ns 0V 136240000.0ns 0V 136280000.0ns 0V 137080000.0ns 0V 137120000.0ns 0V 137520000.0ns 0V 137560000.0ns 0V 138360000.0ns 0V 138400000.0ns 1.95V 138800000.0ns 1.95V 138840000.0ns 0V 139640000.0ns 0V 139680000.0ns 0V 140080000.0ns 0V 140120000.0ns 0V 140920000.0ns 0V 140960000.0ns 0V 141360000.0ns 0V 141400000.0ns 0V 142200000.0ns 0V 142240000.0ns 1.95V 142640000.0ns 1.95V 142680000.0ns 0V 143480000.0ns 0V 143520000.0ns 0V 143920000.0ns 0V 143960000.0ns 0V 144760000.0ns 0V 144800000.0ns 0V 145200000.0ns 0V 145240000.0ns 0V 146040000.0ns 0V 146080000.0ns 1.95V 146480000.0ns 1.95V 146520000.0ns 0V 147320000.0ns 0V 147360000.0ns 0V 147760000.0ns 0V 147800000.0ns 0V 148600000.0ns 0V 148640000.0ns 0V 149040000.0ns 0V 149080000.0ns 0V 149880000.0ns 0V 149920000.0ns 1.95V 150320000.0ns 1.95V 150360000.0ns 0V 151160000.0ns 0V 151200000.0ns 0V 151600000.0ns 0V 151640000.0ns 0V 152440000.0ns 0V 152480000.0ns 0V 152880000.0ns 0V 152920000.0ns 0V 153720000.0ns 0V 153760000.0ns 1.95V 154160000.0ns 1.95V 154200000.0ns 0V 155000000.0ns 0V 155040000.0ns 0V 155440000.0ns 0V 155480000.0ns 0V 156280000.0ns 0V 156320000.0ns 0V 156720000.0ns 0V 156760000.0ns 0V 157560000.0ns 0V 157600000.0ns 1.95V 158000000.0ns 1.95V 158040000.0ns 0V 158840000.0ns 0V 158880000.0ns 0V 159280000.0ns 0V 159320000.0ns 0V 160120000.0ns 0V 160160000.0ns 0V 160560000.0ns 0V 160600000.0ns 0V 161400000.0ns 0V 161440000.0ns 1.95V 161840000.0ns 1.95V 161880000.0ns 0V 162680000.0ns 0V 162720000.0ns 0V 163120000.0ns 0V 163160000.0ns 0V 163960000.0ns 0V 164000000.0ns 0V 164400000.0ns 0V 164440000.0ns 0V 165240000.0ns 0V 165280000.0ns 1.95V 165680000.0ns 1.95V 165720000.0ns 0V 166520000.0ns 0V 166560000.0ns 0V 166960000.0ns 0V 167000000.0ns 0V 167800000.0ns 0V 167840000.0ns 0V 168240000.0ns 0V 168280000.0ns 0V 169080000.0ns 0V 169120000.0ns 1.95V 169520000.0ns 1.95V 169560000.0ns 0V 170360000.0ns 0V 170400000.0ns 0V 170800000.0ns 0V 170840000.0ns 0V 171640000.0ns 0V 171680000.0ns 0V 172080000.0ns 0V 172120000.0ns 0V 172920000.0ns 0V 172960000.0ns 1.95V 173360000.0ns 1.95V 173400000.0ns 0V 174200000.0ns 0V 174240000.0ns 0V 174640000.0ns 0V 174680000.0ns 0V 175480000.0ns 0V 175520000.0ns 0V 175920000.0ns 0V 175960000.0ns 0V 176760000.0ns 0V 176800000.0ns 1.95V 177200000.0ns 1.95V 177240000.0ns 0V 178040000.0ns 0V 178080000.0ns 0V 178480000.0ns 0V 178520000.0ns 0V 179320000.0ns 0V 179360000.0ns 0V 179760000.0ns 0V 179800000.0ns 0V 180600000.0ns 0V 180640000.0ns 1.95V 181040000.0ns 1.95V 181080000.0ns 0V 181880000.0ns 0V 181920000.0ns 0V 182320000.0ns 0V 182360000.0ns 0V 183160000.0ns 0V 183200000.0ns 0V 183600000.0ns 0V 183640000.0ns 0V 184440000.0ns 0V 184480000.0ns 1.95V 184880000.0ns 1.95V 184920000.0ns 0V 185720000.0ns 0V 185760000.0ns 0V 186160000.0ns 0V 186200000.0ns 0V 187000000.0ns 0V 187040000.0ns 0V 187440000.0ns 0V 187480000.0ns 0V 188280000.0ns 0V 188320000.0ns 1.95V 188720000.0ns 1.95V 188760000.0ns 0V 189560000.0ns 0V 189600000.0ns 0V 190000000.0ns 0V 190040000.0ns 0V 190840000.0ns 0V 190880000.0ns 0V 191280000.0ns 0V 191320000.0ns 0V 192120000.0ns 0V 192160000.0ns 1.95V 192560000.0ns 1.95V 192600000.0ns 0V 193400000.0ns 0V 193440000.0ns 0V 193840000.0ns 0V 193880000.0ns 0V 194680000.0ns 0V 194720000.0ns 0V 195120000.0ns 0V 195160000.0ns 0V 195960000.0ns 0V 196000000.0ns 1.95V 196400000.0ns 1.95V 196440000.0ns 0V 197240000.0ns 0V 197280000.0ns 0V 197680000.0ns 0V 197720000.0ns 0V 198520000.0ns 0V 198560000.0ns 0V 198960000.0ns 0V 199000000.0ns 0V 199800000.0ns 0V 199840000.0ns 1.95V 200240000.0ns 1.95V 200280000.0ns 0V 201080000.0ns 0V 201120000.0ns 0V 201520000.0ns 0V 201560000.0ns 0V 202360000.0ns 0V 202400000.0ns 0V 202800000.0ns 0V 202840000.0ns 0V 203640000.0ns 0V 203680000.0ns 1.95V 204080000.0ns 1.95V 204120000.0ns 0V 204920000.0ns 0V 204960000.0ns 0V 205360000.0ns 0V 205400000.0ns 0V 206200000.0ns 0V 206240000.0ns 0V 206640000.0ns 0V 206680000.0ns 0V 207480000.0ns 0V 207520000.0ns 1.95V 207920000.0ns 1.95V 207960000.0ns 0V 208760000.0ns 0V 208800000.0ns 0V 209200000.0ns 0V 209240000.0ns 0V 210040000.0ns 0V 210080000.0ns 0V 210480000.0ns 0V 210520000.0ns 0V 211320000.0ns 0V 211360000.0ns 1.95V 211760000.0ns 1.95V 211800000.0ns 0V 212600000.0ns 0V 212640000.0ns 0V 213040000.0ns 0V 213080000.0ns 0V 213880000.0ns 0V 213920000.0ns 0V 214320000.0ns 0V 214360000.0ns 0V 215160000.0ns 0V 215200000.0ns 1.95V 215600000.0ns 1.95V 215640000.0ns 0V 216440000.0ns 0V 216480000.0ns 0V 216880000.0ns 0V 216920000.0ns 0V 217720000.0ns 0V 217760000.0ns 0V 218160000.0ns 0V 218200000.0ns 0V 219000000.0ns 0V 219040000.0ns 1.95V 219440000.0ns 1.95V 219480000.0ns 0V 220280000.0ns 0V 220320000.0ns 0V 220720000.0ns 0V 220760000.0ns 0V 221560000.0ns 0V 221600000.0ns 0V 222000000.0ns 0V 222040000.0ns 0V 222840000.0ns 0V 222880000.0ns 1.95V 223280000.0ns 1.95V 223320000.0ns 0V 224120000.0ns 0V 224160000.0ns 0V 224560000.0ns 0V 224600000.0ns 0V 225400000.0ns 0V 225440000.0ns 0V 225840000.0ns 0V 225880000.0ns 0V 226680000.0ns 0V 226720000.0ns 1.95V 227120000.0ns 1.95V 227160000.0ns 0V 227960000.0ns 0V 228000000.0ns 0V 228400000.0ns 0V 228440000.0ns 0V 229240000.0ns 0V 229280000.0ns 0V 229680000.0ns 0V 229720000.0ns 0V 230520000.0ns 0V 230560000.0ns 1.95V 230960000.0ns 1.95V 231000000.0ns 0V 231800000.0ns 0V 231840000.0ns 0V 232240000.0ns 0V 232280000.0ns 0V 233080000.0ns 0V 233120000.0ns 0V 233520000.0ns 0V 233560000.0ns 0V 234360000.0ns 0V 234400000.0ns 1.95V 234800000.0ns 1.95V 234840000.0ns 0V 235640000.0ns 0V 235680000.0ns 0V 236080000.0ns 0V 236120000.0ns 0V 236920000.0ns 0V 236960000.0ns 0V 237360000.0ns 0V 237400000.0ns 0V 238200000.0ns 0V 238240000.0ns 1.95V 238640000.0ns 1.95V 238680000.0ns 0V 239480000.0ns 0V 239520000.0ns 0V 239920000.0ns 0V 239960000.0ns 0V 240760000.0ns 0V 240800000.0ns 0V 241200000.0ns 0V 241240000.0ns 0V 242040000.0ns 0V 242080000.0ns 1.95V 242480000.0ns 1.95V 242520000.0ns 0V 243320000.0ns 0V 243360000.0ns 0V 243760000.0ns 0V 243800000.0ns 0V 244600000.0ns 0V 244640000.0ns 0V 245040000.0ns 0V 245080000.0ns 0V 245880000.0ns 0V 245920000.0ns 1.95V 246320000.0ns 1.95V 246360000.0ns 0V 247160000.0ns 0V 247200000.0ns 0V 247600000.0ns 0V 247640000.0ns 0V 248440000.0ns 0V 248480000.0ns 0V 248880000.0ns 0V 248920000.0ns 0V 249720000.0ns 0V 249760000.0ns 1.95V 250160000.0ns 1.95V 250200000.0ns 0V 251000000.0ns 0V 251040000.0ns 0V 251440000.0ns 0V 251480000.0ns 0V 252280000.0ns 0V 252320000.0ns 0V 252720000.0ns 0V 252760000.0ns 0V 253560000.0ns 0V 253600000.0ns 1.95V 254000000.0ns 1.95V 254040000.0ns 0V 254840000.0ns 0V 254880000.0ns 0V 255280000.0ns 0V 255320000.0ns 0V 256120000.0ns 0V 256160000.0ns 0V 256560000.0ns 0V 256600000.0ns 0V 257400000.0ns 0V 257440000.0ns 1.95V 257840000.0ns 1.95V 257880000.0ns 0V 258680000.0ns 0V 258720000.0ns 0V 259120000.0ns 0V 259160000.0ns 0V 259960000.0ns 0V 260000000.0ns 0V 260400000.0ns 0V 260440000.0ns 0V 261240000.0ns 0V 261280000.0ns 1.95V 261680000.0ns 1.95V 261720000.0ns 0V 262520000.0ns 0V 262560000.0ns 0V 262960000.0ns 0V 263000000.0ns 0V 263800000.0ns 0V 263840000.0ns 0V 264240000.0ns 0V 264280000.0ns 0V 265080000.0ns 0V 265120000.0ns 1.95V 265520000.0ns 1.95V 265560000.0ns 0V 266360000.0ns 0V 266400000.0ns 0V 266800000.0ns 0V 266840000.0ns 0V 267640000.0ns 0V 267680000.0ns 0V 268080000.0ns 0V 268120000.0ns 0V 268920000.0ns 0V 268960000.0ns 1.95V 269360000.0ns 1.95V 269400000.0ns 0V 270200000.0ns 0V 270240000.0ns 0V 270640000.0ns 0V 270680000.0ns 0V 271480000.0ns 0V 271520000.0ns 0V 271920000.0ns 0V 271960000.0ns 0V 272760000.0ns 0V 272800000.0ns 1.95V 273200000.0ns 1.95V 273240000.0ns 0V 274040000.0ns 0V 274080000.0ns 0V 274480000.0ns 0V 274520000.0ns 0V 275320000.0ns 0V 275360000.0ns 0V 275760000.0ns 0V 275800000.0ns 0V 276600000.0ns 0V 276640000.0ns 1.95V 277040000.0ns 1.95V 277080000.0ns 0V 277880000.0ns 0V 277920000.0ns 0V 278320000.0ns 0V 278360000.0ns 0V 279160000.0ns 0V 279200000.0ns 0V 279600000.0ns 0V 279640000.0ns 0V 280440000.0ns 0V 280480000.0ns 1.95V 280880000.0ns 1.95V 280920000.0ns 0V 281720000.0ns 0V 281760000.0ns 0V 282160000.0ns 0V 282200000.0ns 0V 283000000.0ns 0V 283040000.0ns 0V 283440000.0ns 0V 283480000.0ns 0V 284280000.0ns 0V 284320000.0ns 1.95V 284720000.0ns 1.95V 284760000.0ns 0V 285560000.0ns 0V 285600000.0ns 0V 286000000.0ns 0V 286040000.0ns 0V 286840000.0ns 0V 286880000.0ns 0V 287280000.0ns 0V 287320000.0ns 0V 288120000.0ns 0V 288160000.0ns 1.95V 288560000.0ns 1.95V 288600000.0ns 0V 289400000.0ns 0V 289440000.0ns 0V 289840000.0ns 0V 289880000.0ns 0V 290680000.0ns 0V 290720000.0ns 0V 291120000.0ns 0V 291160000.0ns 0V 291960000.0ns 0V 292000000.0ns 1.95V 292400000.0ns 1.95V 292440000.0ns 0V 293240000.0ns 0V 293280000.0ns 0V 293680000.0ns 0V 293720000.0ns 0V 294520000.0ns 0V 294560000.0ns 0V 294960000.0ns 0V 295000000.0ns 0V 295800000.0ns 0V 295840000.0ns 1.95V 296240000.0ns 1.95V 296280000.0ns 0V 297080000.0ns 0V 297120000.0ns 0V 297520000.0ns 0V 297560000.0ns 0V 298360000.0ns 0V 298400000.0ns 0V 298800000.0ns 0V 298840000.0ns 0V 299640000.0ns 0V 299680000.0ns 1.95V 300080000.0ns 1.95V 300120000.0ns 0V 300920000.0ns 0V 300960000.0ns 0V 301360000.0ns 0V 301400000.0ns 0V 302200000.0ns 0V 302240000.0ns 0V 302640000.0ns 0V 302680000.0ns 0V 303480000.0ns 0V 303520000.0ns 1.95V 303920000.0ns 1.95V 303960000.0ns 0V 304760000.0ns 0V 304800000.0ns 0V 305200000.0ns 0V 305240000.0ns 0V 306040000.0ns 0V 306080000.0ns 0V 306480000.0ns 0V 306520000.0ns 0V 307320000.0ns 0V 307360000.0ns 1.95V 307760000.0ns 1.95V 307800000.0ns 0V 308600000.0ns 0V 308640000.0ns 0V 309040000.0ns 0V 309080000.0ns 0V 309880000.0ns 0V 309920000.0ns 0V 310320000.0ns 0V 310360000.0ns 0V 311160000.0ns 0V 311200000.0ns 1.95V 311600000.0ns 1.95V 311640000.0ns 0V 312440000.0ns 0V 312480000.0ns 0V 312880000.0ns 0V 312920000.0ns 0V 313720000.0ns 0V 313760000.0ns 0V 314160000.0ns 0V 314200000.0ns 0V 315000000.0ns 0V 315040000.0ns 1.95V 315440000.0ns 1.95V 315480000.0ns 0V 316280000.0ns 0V 316320000.0ns 0V 316720000.0ns 0V 316760000.0ns 0V 317560000.0ns 0V 317600000.0ns 0V 318000000.0ns 0V 318040000.0ns 0V 318840000.0ns 0V 318880000.0ns 1.95V 319280000.0ns 1.95V 319320000.0ns 0V 320120000.0ns 0V 320160000.0ns 0V 320560000.0ns 0V 320600000.0ns 0V 321400000.0ns 0V 321440000.0ns 0V 321840000.0ns 0V 321880000.0ns 0V 322680000.0ns 0V 322720000.0ns 1.95V 323120000.0ns 1.95V 323160000.0ns 0V 323960000.0ns 0V 324000000.0ns 0V 324400000.0ns 0V 324440000.0ns 0V 325240000.0ns 0V 325280000.0ns 0V 325680000.0ns 0V 325720000.0ns 0V 326520000.0ns 0V 326560000.0ns 1.95V 326960000.0ns 1.95V 327000000.0ns 0V 327800000.0ns 0V 327840000.0ns 0V 328240000.0ns 0V 328280000.0ns 0V 329080000.0ns 0V 329120000.0ns 0V 329520000.0ns 0V 329560000.0ns 0V 330360000.0ns 0V 330400000.0ns 1.95V 330800000.0ns 1.95V 330840000.0ns 0V 331640000.0ns 0V 331680000.0ns 0V 332080000.0ns 0V 332120000.0ns 0V 332920000.0ns 0V 332960000.0ns 0V 333360000.0ns 0V 333400000.0ns 0V 334200000.0ns 0V 334240000.0ns 1.95V 334640000.0ns 1.95V 334680000.0ns 0V 335480000.0ns 0V 335520000.0ns 0V 335920000.0ns 0V 335960000.0ns 0V 336760000.0ns 0V 336800000.0ns 0V 337200000.0ns 0V 337240000.0ns 0V 338040000.0ns 0V 338080000.0ns 1.95V 338480000.0ns 1.95V 338520000.0ns 0V 339320000.0ns 0V 339360000.0ns 0V 339760000.0ns 0V 339800000.0ns 0V 340600000.0ns 0V 340640000.0ns 0V 341040000.0ns 0V 341080000.0ns 0V 341880000.0ns 0V 341920000.0ns 1.95V 342320000.0ns 1.95V 342360000.0ns 0V 343160000.0ns 0V 343200000.0ns 0V 343600000.0ns 0V 343640000.0ns 0V 344440000.0ns 0V 344480000.0ns 0V 344880000.0ns 0V 344920000.0ns 0V 345720000.0ns 0V 345760000.0ns 1.95V 346160000.0ns 1.95V 346200000.0ns 0V 347000000.0ns 0V 347040000.0ns 0V 347440000.0ns 0V 347480000.0ns 0V 348280000.0ns 0V 348320000.0ns 0V 348720000.0ns 0V 348760000.0ns 0V 349560000.0ns 0V 349600000.0ns 1.95V 350000000.0ns 1.95V 350040000.0ns 0V 350840000.0ns 0V 350880000.0ns 0V 351280000.0ns 0V 351320000.0ns 0V 352120000.0ns 0V 352160000.0ns 0V 352560000.0ns 0V 352600000.0ns 0V 353400000.0ns 0V 353440000.0ns 1.95V 353840000.0ns 1.95V 353880000.0ns 0V 354680000.0ns 0V 354720000.0ns 0V 355120000.0ns 0V 355160000.0ns 0V 355960000.0ns 0V 356000000.0ns 0V 356400000.0ns 0V 356440000.0ns 0V 357240000.0ns 0V 357280000.0ns 1.95V 357680000.0ns 1.95V 357720000.0ns 0V 358520000.0ns 0V 358560000.0ns 0V 358960000.0ns 0V 359000000.0ns 0V 359800000.0ns 0V 359840000.0ns 0V 360240000.0ns 0V 360280000.0ns 0V 361080000.0ns 0V 361120000.0ns 1.95V 361520000.0ns 1.95V 361560000.0ns 0V 362360000.0ns 0V 362400000.0ns 0V 362800000.0ns 0V 362840000.0ns 0V 363640000.0ns 0V 363680000.0ns 0V 364080000.0ns 0V 364120000.0ns 0V 364920000.0ns 0V 364960000.0ns 1.95V 365360000.0ns 1.95V 365400000.0ns 0V 366200000.0ns 0V 366240000.0ns 0V 366640000.0ns 0V 366680000.0ns 0V 367480000.0ns 0V 367520000.0ns 0V 367920000.0ns 0V 367960000.0ns 0V 368760000.0ns 0V 368800000.0ns 1.95V 369200000.0ns 1.95V 369240000.0ns 0V 370040000.0ns 0V 370080000.0ns 0V 370480000.0ns 0V 370520000.0ns 0V 371320000.0ns 0V 371360000.0ns 0V 371760000.0ns 0V 371800000.0ns 0V 372600000.0ns 0V 372640000.0ns 1.95V 373040000.0ns 1.95V 373080000.0ns 0V 373880000.0ns 0V 373920000.0ns 0V 374320000.0ns 0V 374360000.0ns 0V 375160000.0ns 0V 375200000.0ns 0V 375600000.0ns 0V 375640000.0ns 0V 376440000.0ns 0V 376480000.0ns 1.95V 376880000.0ns 1.95V 376920000.0ns 0V 377720000.0ns 0V 377760000.0ns 0V 378160000.0ns 0V 378200000.0ns 0V 379000000.0ns 0V 379040000.0ns 0V 379440000.0ns 0V 379480000.0ns 0V 380280000.0ns 0V 380320000.0ns 1.95V 380720000.0ns 1.95V 380760000.0ns 0V 381560000.0ns 0V 381600000.0ns 0V 382000000.0ns 0V 382040000.0ns 0V 382840000.0ns 0V 382880000.0ns 0V 383280000.0ns 0V 383320000.0ns 0V 384120000.0ns 0V 384160000.0ns 1.95V 384560000.0ns 1.95V 384600000.0ns 0V 385400000.0ns 0V 385440000.0ns 0V 385840000.0ns 0V 385880000.0ns 0V 386680000.0ns 0V 386720000.0ns 0V 387120000.0ns 0V 387160000.0ns 0V 387960000.0ns 0V 388000000.0ns 1.95V 388400000.0ns 1.95V 388440000.0ns 0V 389240000.0ns 0V 389280000.0ns 0V 389680000.0ns 0V 389720000.0ns 0V 390520000.0ns 0V 390560000.0ns 0V 390960000.0ns 0V 391000000.0ns 0V)
VUPDATE UPDATE 0 PWL(0ns 0V 3960000.0ns 0V 7800000.0ns 0V 7840000.0ns 0V 8240000.0ns 0V 8280000.0ns 0V 9080000.0ns 0V 9120000.0ns 0V 9520000.0ns 0V 9560000.0ns 0V 10360000.0ns 0V 10400000.0ns 1.95V 10800000.0ns 1.95V 10840000.0ns 0V 11640000.0ns 0V 11680000.0ns 0V 12080000.0ns 0V 12120000.0ns 0V 12920000.0ns 0V 12960000.0ns 0V 13360000.0ns 0V 13400000.0ns 0V 14200000.0ns 0V 14240000.0ns 1.95V 14640000.0ns 1.95V 14680000.0ns 0V 15480000.0ns 0V 15520000.0ns 0V 15920000.0ns 0V 15960000.0ns 0V 16760000.0ns 0V 16800000.0ns 0V 17200000.0ns 0V 17240000.0ns 0V 18040000.0ns 0V 18080000.0ns 1.95V 18480000.0ns 1.95V 18520000.0ns 0V 19320000.0ns 0V 19360000.0ns 0V 19760000.0ns 0V 19800000.0ns 0V 20600000.0ns 0V 20640000.0ns 0V 21040000.0ns 0V 21080000.0ns 0V 21880000.0ns 0V 21920000.0ns 1.95V 22320000.0ns 1.95V 22360000.0ns 0V 23160000.0ns 0V 23200000.0ns 0V 23600000.0ns 0V 23640000.0ns 0V 24440000.0ns 0V 24480000.0ns 0V 24880000.0ns 0V 24920000.0ns 0V 25720000.0ns 0V 25760000.0ns 1.95V 26160000.0ns 1.95V 26200000.0ns 0V 27000000.0ns 0V 27040000.0ns 0V 27440000.0ns 0V 27480000.0ns 0V 28280000.0ns 0V 28320000.0ns 0V 28720000.0ns 0V 28760000.0ns 0V 29560000.0ns 0V 29600000.0ns 1.95V 30000000.0ns 1.95V 30040000.0ns 0V 30840000.0ns 0V 30880000.0ns 0V 31280000.0ns 0V 31320000.0ns 0V 32120000.0ns 0V 32160000.0ns 0V 32560000.0ns 0V 32600000.0ns 0V 33400000.0ns 0V 33440000.0ns 1.95V 33840000.0ns 1.95V 33880000.0ns 0V 34680000.0ns 0V 34720000.0ns 0V 35120000.0ns 0V 35160000.0ns 0V 35960000.0ns 0V 36000000.0ns 0V 36400000.0ns 0V 36440000.0ns 0V 37240000.0ns 0V 37280000.0ns 1.95V 37680000.0ns 1.95V 37720000.0ns 0V 38520000.0ns 0V 38560000.0ns 0V 38960000.0ns 0V 39000000.0ns 0V 39800000.0ns 0V 39840000.0ns 0V 40240000.0ns 0V 40280000.0ns 0V 41080000.0ns 0V 41120000.0ns 1.95V 41520000.0ns 1.95V 41560000.0ns 0V 42360000.0ns 0V 42400000.0ns 0V 42800000.0ns 0V 42840000.0ns 0V 43640000.0ns 0V 43680000.0ns 0V 44080000.0ns 0V 44120000.0ns 0V 44920000.0ns 0V 44960000.0ns 1.95V 45360000.0ns 1.95V 45400000.0ns 0V 46200000.0ns 0V 46240000.0ns 0V 46640000.0ns 0V 46680000.0ns 0V 47480000.0ns 0V 47520000.0ns 0V 47920000.0ns 0V 47960000.0ns 0V 48760000.0ns 0V 48800000.0ns 1.95V 49200000.0ns 1.95V 49240000.0ns 0V 50040000.0ns 0V 50080000.0ns 0V 50480000.0ns 0V 50520000.0ns 0V 51320000.0ns 0V 51360000.0ns 0V 51760000.0ns 0V 51800000.0ns 0V 52600000.0ns 0V 52640000.0ns 1.95V 53040000.0ns 1.95V 53080000.0ns 0V 53880000.0ns 0V 53920000.0ns 0V 54320000.0ns 0V 54360000.0ns 0V 55160000.0ns 0V 55200000.0ns 0V 55600000.0ns 0V 55640000.0ns 0V 56440000.0ns 0V 56480000.0ns 1.95V 56880000.0ns 1.95V 56920000.0ns 0V 57720000.0ns 0V 57760000.0ns 0V 58160000.0ns 0V 58200000.0ns 0V 59000000.0ns 0V 59040000.0ns 0V 59440000.0ns 0V 59480000.0ns 0V 60280000.0ns 0V 60320000.0ns 1.95V 60720000.0ns 1.95V 60760000.0ns 0V 61560000.0ns 0V 61600000.0ns 0V 62000000.0ns 0V 62040000.0ns 0V 62840000.0ns 0V 62880000.0ns 0V 63280000.0ns 0V 63320000.0ns 0V 64120000.0ns 0V 64160000.0ns 1.95V 64560000.0ns 1.95V 64600000.0ns 0V 65400000.0ns 0V 65440000.0ns 0V 65840000.0ns 0V 65880000.0ns 0V 66680000.0ns 0V 66720000.0ns 0V 67120000.0ns 0V 67160000.0ns 0V 67960000.0ns 0V 68000000.0ns 1.95V 68400000.0ns 1.95V 68440000.0ns 0V 69240000.0ns 0V 69280000.0ns 0V 69680000.0ns 0V 69720000.0ns 0V 70520000.0ns 0V 70560000.0ns 0V 70960000.0ns 0V 71000000.0ns 0V 71800000.0ns 0V 71840000.0ns 1.95V 72240000.0ns 1.95V 72280000.0ns 0V 73080000.0ns 0V 73120000.0ns 0V 73520000.0ns 0V 73560000.0ns 0V 74360000.0ns 0V 74400000.0ns 0V 74800000.0ns 0V 74840000.0ns 0V 75640000.0ns 0V 75680000.0ns 1.95V 76080000.0ns 1.95V 76120000.0ns 0V 76920000.0ns 0V 76960000.0ns 0V 77360000.0ns 0V 77400000.0ns 0V 78200000.0ns 0V 78240000.0ns 0V 78640000.0ns 0V 78680000.0ns 0V 79480000.0ns 0V 79520000.0ns 1.95V 79920000.0ns 1.95V 79960000.0ns 0V 80760000.0ns 0V 80800000.0ns 0V 81200000.0ns 0V 81240000.0ns 0V 82040000.0ns 0V 82080000.0ns 0V 82480000.0ns 0V 82520000.0ns 0V 83320000.0ns 0V 83360000.0ns 1.95V 83760000.0ns 1.95V 83800000.0ns 0V 84600000.0ns 0V 84640000.0ns 0V 85040000.0ns 0V 85080000.0ns 0V 85880000.0ns 0V 85920000.0ns 0V 86320000.0ns 0V 86360000.0ns 0V 87160000.0ns 0V 87200000.0ns 1.95V 87600000.0ns 1.95V 87640000.0ns 0V 88440000.0ns 0V 88480000.0ns 0V 88880000.0ns 0V 88920000.0ns 0V 89720000.0ns 0V 89760000.0ns 0V 90160000.0ns 0V 90200000.0ns 0V 91000000.0ns 0V 91040000.0ns 1.95V 91440000.0ns 1.95V 91480000.0ns 0V 92280000.0ns 0V 92320000.0ns 0V 92720000.0ns 0V 92760000.0ns 0V 93560000.0ns 0V 93600000.0ns 0V 94000000.0ns 0V 94040000.0ns 0V 94840000.0ns 0V 94880000.0ns 1.95V 95280000.0ns 1.95V 95320000.0ns 0V 96120000.0ns 0V 96160000.0ns 0V 96560000.0ns 0V 96600000.0ns 0V 97400000.0ns 0V 97440000.0ns 0V 97840000.0ns 0V 97880000.0ns 0V 98680000.0ns 0V 98720000.0ns 1.95V 99120000.0ns 1.95V 99160000.0ns 0V 99960000.0ns 0V 100000000.0ns 0V 100400000.0ns 0V 100440000.0ns 0V 101240000.0ns 0V 101280000.0ns 0V 101680000.0ns 0V 101720000.0ns 0V 102520000.0ns 0V 102560000.0ns 1.95V 102960000.0ns 1.95V 103000000.0ns 0V 103800000.0ns 0V 103840000.0ns 0V 104240000.0ns 0V 104280000.0ns 0V 105080000.0ns 0V 105120000.0ns 0V 105520000.0ns 0V 105560000.0ns 0V 106360000.0ns 0V 106400000.0ns 1.95V 106800000.0ns 1.95V 106840000.0ns 0V 107640000.0ns 0V 107680000.0ns 0V 108080000.0ns 0V 108120000.0ns 0V 108920000.0ns 0V 108960000.0ns 0V 109360000.0ns 0V 109400000.0ns 0V 110200000.0ns 0V 110240000.0ns 1.95V 110640000.0ns 1.95V 110680000.0ns 0V 111480000.0ns 0V 111520000.0ns 0V 111920000.0ns 0V 111960000.0ns 0V 112760000.0ns 0V 112800000.0ns 0V 113200000.0ns 0V 113240000.0ns 0V 114040000.0ns 0V 114080000.0ns 1.95V 114480000.0ns 1.95V 114520000.0ns 0V 115320000.0ns 0V 115360000.0ns 0V 115760000.0ns 0V 115800000.0ns 0V 116600000.0ns 0V 116640000.0ns 0V 117040000.0ns 0V 117080000.0ns 0V 117880000.0ns 0V 117920000.0ns 1.95V 118320000.0ns 1.95V 118360000.0ns 0V 119160000.0ns 0V 119200000.0ns 0V 119600000.0ns 0V 119640000.0ns 0V 120440000.0ns 0V 120480000.0ns 0V 120880000.0ns 0V 120920000.0ns 0V 121720000.0ns 0V 121760000.0ns 1.95V 122160000.0ns 1.95V 122200000.0ns 0V 123000000.0ns 0V 123040000.0ns 0V 123440000.0ns 0V 123480000.0ns 0V 124280000.0ns 0V 124320000.0ns 0V 124720000.0ns 0V 124760000.0ns 0V 125560000.0ns 0V 125600000.0ns 1.95V 126000000.0ns 1.95V 126040000.0ns 0V 126840000.0ns 0V 126880000.0ns 0V 127280000.0ns 0V 127320000.0ns 0V 128120000.0ns 0V 128160000.0ns 0V 128560000.0ns 0V 128600000.0ns 0V 129400000.0ns 0V 129440000.0ns 1.95V 129840000.0ns 1.95V 129880000.0ns 0V 130680000.0ns 0V 130720000.0ns 0V 131120000.0ns 0V 131160000.0ns 0V 131960000.0ns 0V 132000000.0ns 0V 132400000.0ns 0V 132440000.0ns 0V 133240000.0ns 0V 133280000.0ns 1.95V 133680000.0ns 1.95V 133720000.0ns 0V 134520000.0ns 0V 134560000.0ns 0V 134960000.0ns 0V 135000000.0ns 0V 135800000.0ns 0V 135840000.0ns 0V 136240000.0ns 0V 136280000.0ns 0V 137080000.0ns 0V 137120000.0ns 1.95V 137520000.0ns 1.95V 137560000.0ns 0V 138360000.0ns 0V 138400000.0ns 0V 138800000.0ns 0V 138840000.0ns 0V 139640000.0ns 0V 139680000.0ns 0V 140080000.0ns 0V 140120000.0ns 0V 140920000.0ns 0V 140960000.0ns 1.95V 141360000.0ns 1.95V 141400000.0ns 0V 142200000.0ns 0V 142240000.0ns 0V 142640000.0ns 0V 142680000.0ns 0V 143480000.0ns 0V 143520000.0ns 0V 143920000.0ns 0V 143960000.0ns 0V 144760000.0ns 0V 144800000.0ns 1.95V 145200000.0ns 1.95V 145240000.0ns 0V 146040000.0ns 0V 146080000.0ns 0V 146480000.0ns 0V 146520000.0ns 0V 147320000.0ns 0V 147360000.0ns 0V 147760000.0ns 0V 147800000.0ns 0V 148600000.0ns 0V 148640000.0ns 1.95V 149040000.0ns 1.95V 149080000.0ns 0V 149880000.0ns 0V 149920000.0ns 0V 150320000.0ns 0V 150360000.0ns 0V 151160000.0ns 0V 151200000.0ns 0V 151600000.0ns 0V 151640000.0ns 0V 152440000.0ns 0V 152480000.0ns 1.95V 152880000.0ns 1.95V 152920000.0ns 0V 153720000.0ns 0V 153760000.0ns 0V 154160000.0ns 0V 154200000.0ns 0V 155000000.0ns 0V 155040000.0ns 0V 155440000.0ns 0V 155480000.0ns 0V 156280000.0ns 0V 156320000.0ns 1.95V 156720000.0ns 1.95V 156760000.0ns 0V 157560000.0ns 0V 157600000.0ns 0V 158000000.0ns 0V 158040000.0ns 0V 158840000.0ns 0V 158880000.0ns 0V 159280000.0ns 0V 159320000.0ns 0V 160120000.0ns 0V 160160000.0ns 1.95V 160560000.0ns 1.95V 160600000.0ns 0V 161400000.0ns 0V 161440000.0ns 0V 161840000.0ns 0V 161880000.0ns 0V 162680000.0ns 0V 162720000.0ns 0V 163120000.0ns 0V 163160000.0ns 0V 163960000.0ns 0V 164000000.0ns 1.95V 164400000.0ns 1.95V 164440000.0ns 0V 165240000.0ns 0V 165280000.0ns 0V 165680000.0ns 0V 165720000.0ns 0V 166520000.0ns 0V 166560000.0ns 0V 166960000.0ns 0V 167000000.0ns 0V 167800000.0ns 0V 167840000.0ns 1.95V 168240000.0ns 1.95V 168280000.0ns 0V 169080000.0ns 0V 169120000.0ns 0V 169520000.0ns 0V 169560000.0ns 0V 170360000.0ns 0V 170400000.0ns 0V 170800000.0ns 0V 170840000.0ns 0V 171640000.0ns 0V 171680000.0ns 1.95V 172080000.0ns 1.95V 172120000.0ns 0V 172920000.0ns 0V 172960000.0ns 0V 173360000.0ns 0V 173400000.0ns 0V 174200000.0ns 0V 174240000.0ns 0V 174640000.0ns 0V 174680000.0ns 0V 175480000.0ns 0V 175520000.0ns 1.95V 175920000.0ns 1.95V 175960000.0ns 0V 176760000.0ns 0V 176800000.0ns 0V 177200000.0ns 0V 177240000.0ns 0V 178040000.0ns 0V 178080000.0ns 0V 178480000.0ns 0V 178520000.0ns 0V 179320000.0ns 0V 179360000.0ns 1.95V 179760000.0ns 1.95V 179800000.0ns 0V 180600000.0ns 0V 180640000.0ns 0V 181040000.0ns 0V 181080000.0ns 0V 181880000.0ns 0V 181920000.0ns 0V 182320000.0ns 0V 182360000.0ns 0V 183160000.0ns 0V 183200000.0ns 1.95V 183600000.0ns 1.95V 183640000.0ns 0V 184440000.0ns 0V 184480000.0ns 0V 184880000.0ns 0V 184920000.0ns 0V 185720000.0ns 0V 185760000.0ns 0V 186160000.0ns 0V 186200000.0ns 0V 187000000.0ns 0V 187040000.0ns 1.95V 187440000.0ns 1.95V 187480000.0ns 0V 188280000.0ns 0V 188320000.0ns 0V 188720000.0ns 0V 188760000.0ns 0V 189560000.0ns 0V 189600000.0ns 0V 190000000.0ns 0V 190040000.0ns 0V 190840000.0ns 0V 190880000.0ns 1.95V 191280000.0ns 1.95V 191320000.0ns 0V 192120000.0ns 0V 192160000.0ns 0V 192560000.0ns 0V 192600000.0ns 0V 193400000.0ns 0V 193440000.0ns 0V 193840000.0ns 0V 193880000.0ns 0V 194680000.0ns 0V 194720000.0ns 1.95V 195120000.0ns 1.95V 195160000.0ns 0V 195960000.0ns 0V 196000000.0ns 0V 196400000.0ns 0V 196440000.0ns 0V 197240000.0ns 0V 197280000.0ns 0V 197680000.0ns 0V 197720000.0ns 0V 198520000.0ns 0V 198560000.0ns 1.95V 198960000.0ns 1.95V 199000000.0ns 0V 199800000.0ns 0V 199840000.0ns 0V 200240000.0ns 0V 200280000.0ns 0V 201080000.0ns 0V 201120000.0ns 0V 201520000.0ns 0V 201560000.0ns 0V 202360000.0ns 0V 202400000.0ns 1.95V 202800000.0ns 1.95V 202840000.0ns 0V 203640000.0ns 0V 203680000.0ns 0V 204080000.0ns 0V 204120000.0ns 0V 204920000.0ns 0V 204960000.0ns 0V 205360000.0ns 0V 205400000.0ns 0V 206200000.0ns 0V 206240000.0ns 1.95V 206640000.0ns 1.95V 206680000.0ns 0V 207480000.0ns 0V 207520000.0ns 0V 207920000.0ns 0V 207960000.0ns 0V 208760000.0ns 0V 208800000.0ns 0V 209200000.0ns 0V 209240000.0ns 0V 210040000.0ns 0V 210080000.0ns 1.95V 210480000.0ns 1.95V 210520000.0ns 0V 211320000.0ns 0V 211360000.0ns 0V 211760000.0ns 0V 211800000.0ns 0V 212600000.0ns 0V 212640000.0ns 0V 213040000.0ns 0V 213080000.0ns 0V 213880000.0ns 0V 213920000.0ns 1.95V 214320000.0ns 1.95V 214360000.0ns 0V 215160000.0ns 0V 215200000.0ns 0V 215600000.0ns 0V 215640000.0ns 0V 216440000.0ns 0V 216480000.0ns 0V 216880000.0ns 0V 216920000.0ns 0V 217720000.0ns 0V 217760000.0ns 1.95V 218160000.0ns 1.95V 218200000.0ns 0V 219000000.0ns 0V 219040000.0ns 0V 219440000.0ns 0V 219480000.0ns 0V 220280000.0ns 0V 220320000.0ns 0V 220720000.0ns 0V 220760000.0ns 0V 221560000.0ns 0V 221600000.0ns 1.95V 222000000.0ns 1.95V 222040000.0ns 0V 222840000.0ns 0V 222880000.0ns 0V 223280000.0ns 0V 223320000.0ns 0V 224120000.0ns 0V 224160000.0ns 0V 224560000.0ns 0V 224600000.0ns 0V 225400000.0ns 0V 225440000.0ns 1.95V 225840000.0ns 1.95V 225880000.0ns 0V 226680000.0ns 0V 226720000.0ns 0V 227120000.0ns 0V 227160000.0ns 0V 227960000.0ns 0V 228000000.0ns 0V 228400000.0ns 0V 228440000.0ns 0V 229240000.0ns 0V 229280000.0ns 1.95V 229680000.0ns 1.95V 229720000.0ns 0V 230520000.0ns 0V 230560000.0ns 0V 230960000.0ns 0V 231000000.0ns 0V 231800000.0ns 0V 231840000.0ns 0V 232240000.0ns 0V 232280000.0ns 0V 233080000.0ns 0V 233120000.0ns 1.95V 233520000.0ns 1.95V 233560000.0ns 0V 234360000.0ns 0V 234400000.0ns 0V 234800000.0ns 0V 234840000.0ns 0V 235640000.0ns 0V 235680000.0ns 0V 236080000.0ns 0V 236120000.0ns 0V 236920000.0ns 0V 236960000.0ns 1.95V 237360000.0ns 1.95V 237400000.0ns 0V 238200000.0ns 0V 238240000.0ns 0V 238640000.0ns 0V 238680000.0ns 0V 239480000.0ns 0V 239520000.0ns 0V 239920000.0ns 0V 239960000.0ns 0V 240760000.0ns 0V 240800000.0ns 1.95V 241200000.0ns 1.95V 241240000.0ns 0V 242040000.0ns 0V 242080000.0ns 0V 242480000.0ns 0V 242520000.0ns 0V 243320000.0ns 0V 243360000.0ns 0V 243760000.0ns 0V 243800000.0ns 0V 244600000.0ns 0V 244640000.0ns 1.95V 245040000.0ns 1.95V 245080000.0ns 0V 245880000.0ns 0V 245920000.0ns 0V 246320000.0ns 0V 246360000.0ns 0V 247160000.0ns 0V 247200000.0ns 0V 247600000.0ns 0V 247640000.0ns 0V 248440000.0ns 0V 248480000.0ns 1.95V 248880000.0ns 1.95V 248920000.0ns 0V 249720000.0ns 0V 249760000.0ns 0V 250160000.0ns 0V 250200000.0ns 0V 251000000.0ns 0V 251040000.0ns 0V 251440000.0ns 0V 251480000.0ns 0V 252280000.0ns 0V 252320000.0ns 1.95V 252720000.0ns 1.95V 252760000.0ns 0V 253560000.0ns 0V 253600000.0ns 0V 254000000.0ns 0V 254040000.0ns 0V 254840000.0ns 0V 254880000.0ns 0V 255280000.0ns 0V 255320000.0ns 0V 256120000.0ns 0V 256160000.0ns 1.95V 256560000.0ns 1.95V 256600000.0ns 0V 257400000.0ns 0V 257440000.0ns 0V 257840000.0ns 0V 257880000.0ns 0V 258680000.0ns 0V 258720000.0ns 0V 259120000.0ns 0V 259160000.0ns 0V 259960000.0ns 0V 260000000.0ns 1.95V 260400000.0ns 1.95V 260440000.0ns 0V 261240000.0ns 0V 261280000.0ns 0V 261680000.0ns 0V 261720000.0ns 0V 262520000.0ns 0V 262560000.0ns 0V 262960000.0ns 0V 263000000.0ns 0V 263800000.0ns 0V 263840000.0ns 1.95V 264240000.0ns 1.95V 264280000.0ns 0V 265080000.0ns 0V 265120000.0ns 0V 265520000.0ns 0V 265560000.0ns 0V 266360000.0ns 0V 266400000.0ns 0V 266800000.0ns 0V 266840000.0ns 0V 267640000.0ns 0V 267680000.0ns 1.95V 268080000.0ns 1.95V 268120000.0ns 0V 268920000.0ns 0V 268960000.0ns 0V 269360000.0ns 0V 269400000.0ns 0V 270200000.0ns 0V 270240000.0ns 0V 270640000.0ns 0V 270680000.0ns 0V 271480000.0ns 0V 271520000.0ns 1.95V 271920000.0ns 1.95V 271960000.0ns 0V 272760000.0ns 0V 272800000.0ns 0V 273200000.0ns 0V 273240000.0ns 0V 274040000.0ns 0V 274080000.0ns 0V 274480000.0ns 0V 274520000.0ns 0V 275320000.0ns 0V 275360000.0ns 1.95V 275760000.0ns 1.95V 275800000.0ns 0V 276600000.0ns 0V 276640000.0ns 0V 277040000.0ns 0V 277080000.0ns 0V 277880000.0ns 0V 277920000.0ns 0V 278320000.0ns 0V 278360000.0ns 0V 279160000.0ns 0V 279200000.0ns 1.95V 279600000.0ns 1.95V 279640000.0ns 0V 280440000.0ns 0V 280480000.0ns 0V 280880000.0ns 0V 280920000.0ns 0V 281720000.0ns 0V 281760000.0ns 0V 282160000.0ns 0V 282200000.0ns 0V 283000000.0ns 0V 283040000.0ns 1.95V 283440000.0ns 1.95V 283480000.0ns 0V 284280000.0ns 0V 284320000.0ns 0V 284720000.0ns 0V 284760000.0ns 0V 285560000.0ns 0V 285600000.0ns 0V 286000000.0ns 0V 286040000.0ns 0V 286840000.0ns 0V 286880000.0ns 1.95V 287280000.0ns 1.95V 287320000.0ns 0V 288120000.0ns 0V 288160000.0ns 0V 288560000.0ns 0V 288600000.0ns 0V 289400000.0ns 0V 289440000.0ns 0V 289840000.0ns 0V 289880000.0ns 0V 290680000.0ns 0V 290720000.0ns 1.95V 291120000.0ns 1.95V 291160000.0ns 0V 291960000.0ns 0V 292000000.0ns 0V 292400000.0ns 0V 292440000.0ns 0V 293240000.0ns 0V 293280000.0ns 0V 293680000.0ns 0V 293720000.0ns 0V 294520000.0ns 0V 294560000.0ns 1.95V 294960000.0ns 1.95V 295000000.0ns 0V 295800000.0ns 0V 295840000.0ns 0V 296240000.0ns 0V 296280000.0ns 0V 297080000.0ns 0V 297120000.0ns 0V 297520000.0ns 0V 297560000.0ns 0V 298360000.0ns 0V 298400000.0ns 1.95V 298800000.0ns 1.95V 298840000.0ns 0V 299640000.0ns 0V 299680000.0ns 0V 300080000.0ns 0V 300120000.0ns 0V 300920000.0ns 0V 300960000.0ns 0V 301360000.0ns 0V 301400000.0ns 0V 302200000.0ns 0V 302240000.0ns 1.95V 302640000.0ns 1.95V 302680000.0ns 0V 303480000.0ns 0V 303520000.0ns 0V 303920000.0ns 0V 303960000.0ns 0V 304760000.0ns 0V 304800000.0ns 0V 305200000.0ns 0V 305240000.0ns 0V 306040000.0ns 0V 306080000.0ns 1.95V 306480000.0ns 1.95V 306520000.0ns 0V 307320000.0ns 0V 307360000.0ns 0V 307760000.0ns 0V 307800000.0ns 0V 308600000.0ns 0V 308640000.0ns 0V 309040000.0ns 0V 309080000.0ns 0V 309880000.0ns 0V 309920000.0ns 1.95V 310320000.0ns 1.95V 310360000.0ns 0V 311160000.0ns 0V 311200000.0ns 0V 311600000.0ns 0V 311640000.0ns 0V 312440000.0ns 0V 312480000.0ns 0V 312880000.0ns 0V 312920000.0ns 0V 313720000.0ns 0V 313760000.0ns 1.95V 314160000.0ns 1.95V 314200000.0ns 0V 315000000.0ns 0V 315040000.0ns 0V 315440000.0ns 0V 315480000.0ns 0V 316280000.0ns 0V 316320000.0ns 0V 316720000.0ns 0V 316760000.0ns 0V 317560000.0ns 0V 317600000.0ns 1.95V 318000000.0ns 1.95V 318040000.0ns 0V 318840000.0ns 0V 318880000.0ns 0V 319280000.0ns 0V 319320000.0ns 0V 320120000.0ns 0V 320160000.0ns 0V 320560000.0ns 0V 320600000.0ns 0V 321400000.0ns 0V 321440000.0ns 1.95V 321840000.0ns 1.95V 321880000.0ns 0V 322680000.0ns 0V 322720000.0ns 0V 323120000.0ns 0V 323160000.0ns 0V 323960000.0ns 0V 324000000.0ns 0V 324400000.0ns 0V 324440000.0ns 0V 325240000.0ns 0V 325280000.0ns 1.95V 325680000.0ns 1.95V 325720000.0ns 0V 326520000.0ns 0V 326560000.0ns 0V 326960000.0ns 0V 327000000.0ns 0V 327800000.0ns 0V 327840000.0ns 0V 328240000.0ns 0V 328280000.0ns 0V 329080000.0ns 0V 329120000.0ns 1.95V 329520000.0ns 1.95V 329560000.0ns 0V 330360000.0ns 0V 330400000.0ns 0V 330800000.0ns 0V 330840000.0ns 0V 331640000.0ns 0V 331680000.0ns 0V 332080000.0ns 0V 332120000.0ns 0V 332920000.0ns 0V 332960000.0ns 1.95V 333360000.0ns 1.95V 333400000.0ns 0V 334200000.0ns 0V 334240000.0ns 0V 334640000.0ns 0V 334680000.0ns 0V 335480000.0ns 0V 335520000.0ns 0V 335920000.0ns 0V 335960000.0ns 0V 336760000.0ns 0V 336800000.0ns 1.95V 337200000.0ns 1.95V 337240000.0ns 0V 338040000.0ns 0V 338080000.0ns 0V 338480000.0ns 0V 338520000.0ns 0V 339320000.0ns 0V 339360000.0ns 0V 339760000.0ns 0V 339800000.0ns 0V 340600000.0ns 0V 340640000.0ns 1.95V 341040000.0ns 1.95V 341080000.0ns 0V 341880000.0ns 0V 341920000.0ns 0V 342320000.0ns 0V 342360000.0ns 0V 343160000.0ns 0V 343200000.0ns 0V 343600000.0ns 0V 343640000.0ns 0V 344440000.0ns 0V 344480000.0ns 1.95V 344880000.0ns 1.95V 344920000.0ns 0V 345720000.0ns 0V 345760000.0ns 0V 346160000.0ns 0V 346200000.0ns 0V 347000000.0ns 0V 347040000.0ns 0V 347440000.0ns 0V 347480000.0ns 0V 348280000.0ns 0V 348320000.0ns 1.95V 348720000.0ns 1.95V 348760000.0ns 0V 349560000.0ns 0V 349600000.0ns 0V 350000000.0ns 0V 350040000.0ns 0V 350840000.0ns 0V 350880000.0ns 0V 351280000.0ns 0V 351320000.0ns 0V 352120000.0ns 0V 352160000.0ns 1.95V 352560000.0ns 1.95V 352600000.0ns 0V 353400000.0ns 0V 353440000.0ns 0V 353840000.0ns 0V 353880000.0ns 0V 354680000.0ns 0V 354720000.0ns 0V 355120000.0ns 0V 355160000.0ns 0V 355960000.0ns 0V 356000000.0ns 1.95V 356400000.0ns 1.95V 356440000.0ns 0V 357240000.0ns 0V 357280000.0ns 0V 357680000.0ns 0V 357720000.0ns 0V 358520000.0ns 0V 358560000.0ns 0V 358960000.0ns 0V 359000000.0ns 0V 359800000.0ns 0V 359840000.0ns 1.95V 360240000.0ns 1.95V 360280000.0ns 0V 361080000.0ns 0V 361120000.0ns 0V 361520000.0ns 0V 361560000.0ns 0V 362360000.0ns 0V 362400000.0ns 0V 362800000.0ns 0V 362840000.0ns 0V 363640000.0ns 0V 363680000.0ns 1.95V 364080000.0ns 1.95V 364120000.0ns 0V 364920000.0ns 0V 364960000.0ns 0V 365360000.0ns 0V 365400000.0ns 0V 366200000.0ns 0V 366240000.0ns 0V 366640000.0ns 0V 366680000.0ns 0V 367480000.0ns 0V 367520000.0ns 1.95V 367920000.0ns 1.95V 367960000.0ns 0V 368760000.0ns 0V 368800000.0ns 0V 369200000.0ns 0V 369240000.0ns 0V 370040000.0ns 0V 370080000.0ns 0V 370480000.0ns 0V 370520000.0ns 0V 371320000.0ns 0V 371360000.0ns 1.95V 371760000.0ns 1.95V 371800000.0ns 0V 372600000.0ns 0V 372640000.0ns 0V 373040000.0ns 0V 373080000.0ns 0V 373880000.0ns 0V 373920000.0ns 0V 374320000.0ns 0V 374360000.0ns 0V 375160000.0ns 0V 375200000.0ns 1.95V 375600000.0ns 1.95V 375640000.0ns 0V 376440000.0ns 0V 376480000.0ns 0V 376880000.0ns 0V 376920000.0ns 0V 377720000.0ns 0V 377760000.0ns 0V 378160000.0ns 0V 378200000.0ns 0V 379000000.0ns 0V 379040000.0ns 1.95V 379440000.0ns 1.95V 379480000.0ns 0V 380280000.0ns 0V 380320000.0ns 0V 380720000.0ns 0V 380760000.0ns 0V 381560000.0ns 0V 381600000.0ns 0V 382000000.0ns 0V 382040000.0ns 0V 382840000.0ns 0V 382880000.0ns 1.95V 383280000.0ns 1.95V 383320000.0ns 0V 384120000.0ns 0V 384160000.0ns 0V 384560000.0ns 0V 384600000.0ns 0V 385400000.0ns 0V 385440000.0ns 0V 385840000.0ns 0V 385880000.0ns 0V 386680000.0ns 0V 386720000.0ns 1.95V 387120000.0ns 1.95V 387160000.0ns 0V 387960000.0ns 0V 388000000.0ns 0V 388400000.0ns 0V 388440000.0ns 0V 389240000.0ns 0V 389280000.0ns 0V 389680000.0ns 0V 389720000.0ns 0V 390520000.0ns 0V 390560000.0ns 1.95V 390960000.0ns 1.95V 391000000.0ns 0V)
VX_0 X_0 0 PWL(0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0.18092870712280273V 8400000.0ns 0.18092870712280273V 8440000.0ns 0.18092870712280273V 8920000.0ns 0.18092870712280273V 8960000.0ns 0.18092870712280273V 9680000.0ns 0.18092870712280273V 9720000.0ns 0.18092870712280273V 10200000.0ns 0.18092870712280273V 10240000.0ns 0.18092870712280273V 10960000.0ns 0.18092870712280273V 11000000.0ns 0V 11480000.0ns 0V 11520000.0ns 0.3246403932571411V 12240000.0ns 0.3246403932571411V 12280000.0ns 0.3246403932571411V 12760000.0ns 0.3246403932571411V 12800000.0ns 0.3246403932571411V 13520000.0ns 0.3246403932571411V 13560000.0ns 0.3246403932571411V 14040000.0ns 0.3246403932571411V 14080000.0ns 0.3246403932571411V 14800000.0ns 0.3246403932571411V 14840000.0ns 0V 15320000.0ns 0V 15360000.0ns 1.9728596210479736V 16080000.0ns 1.9728596210479736V 16120000.0ns 1.9728596210479736V 16600000.0ns 1.9728596210479736V 16640000.0ns 1.9728596210479736V 17360000.0ns 1.9728596210479736V 17400000.0ns 1.9728596210479736V 17880000.0ns 1.9728596210479736V 17920000.0ns 1.9728596210479736V 18640000.0ns 1.9728596210479736V 18680000.0ns 0V 19160000.0ns 0V 19200000.0ns 0.9325268268585205V 19920000.0ns 0.9325268268585205V 19960000.0ns 0.9325268268585205V 20440000.0ns 0.9325268268585205V 20480000.0ns 0.9325268268585205V 21200000.0ns 0.9325268268585205V 21240000.0ns 0.9325268268585205V 21720000.0ns 0.9325268268585205V 21760000.0ns 0.9325268268585205V 22480000.0ns 0.9325268268585205V 22520000.0ns 0V 23000000.0ns 0V 23040000.0ns 0.38829612731933594V 23760000.0ns 0.38829612731933594V 23800000.0ns 0.38829612731933594V 24280000.0ns 0.38829612731933594V 24320000.0ns 0.38829612731933594V 25040000.0ns 0.38829612731933594V 25080000.0ns 0.38829612731933594V 25560000.0ns 0.38829612731933594V 25600000.0ns 0.38829612731933594V 26320000.0ns 0.38829612731933594V 26360000.0ns 0V 26840000.0ns 0V 26880000.0ns 1.8211740255355835V 27600000.0ns 1.8211740255355835V 27640000.0ns 1.8211740255355835V 28120000.0ns 1.8211740255355835V 28160000.0ns 1.8211740255355835V 28880000.0ns 1.8211740255355835V 28920000.0ns 1.8211740255355835V 29400000.0ns 1.8211740255355835V 29440000.0ns 1.8211740255355835V 30160000.0ns 1.8211740255355835V 30200000.0ns 0V 30680000.0ns 0V 30720000.0ns 1.3780229091644287V 31440000.0ns 1.3780229091644287V 31480000.0ns 1.3780229091644287V 31960000.0ns 1.3780229091644287V 32000000.0ns 1.3780229091644287V 32720000.0ns 1.3780229091644287V 32760000.0ns 1.3780229091644287V 33240000.0ns 1.3780229091644287V 33280000.0ns 1.3780229091644287V 34000000.0ns 1.3780229091644287V 34040000.0ns 0V 34520000.0ns 0V 34560000.0ns 1.9736623764038086V 35280000.0ns 1.9736623764038086V 35320000.0ns 1.9736623764038086V 35800000.0ns 1.9736623764038086V 35840000.0ns 1.9736623764038086V 36560000.0ns 1.9736623764038086V 36600000.0ns 1.9736623764038086V 37080000.0ns 1.9736623764038086V 37120000.0ns 1.9736623764038086V 37840000.0ns 1.9736623764038086V 37880000.0ns 0V 38360000.0ns 0V 38400000.0ns 0.06996047496795654V 39120000.0ns 0.06996047496795654V 39160000.0ns 0.06996047496795654V 39640000.0ns 0.06996047496795654V 39680000.0ns 0.06996047496795654V 40400000.0ns 0.06996047496795654V 40440000.0ns 0.06996047496795654V 40920000.0ns 0.06996047496795654V 40960000.0ns 0.06996047496795654V 41680000.0ns 0.06996047496795654V 41720000.0ns 0V 42200000.0ns 0V 42240000.0ns 0.4799463748931885V 42960000.0ns 0.4799463748931885V 43000000.0ns 0.4799463748931885V 43480000.0ns 0.4799463748931885V 43520000.0ns 0.4799463748931885V 44240000.0ns 0.4799463748931885V 44280000.0ns 0.4799463748931885V 44760000.0ns 0.4799463748931885V 44800000.0ns 0.4799463748931885V 45520000.0ns 0.4799463748931885V 45560000.0ns 0V 46040000.0ns 0V 46080000.0ns 0.20705318450927734V 46800000.0ns 0.20705318450927734V 46840000.0ns 0.20705318450927734V 47320000.0ns 0.20705318450927734V 47360000.0ns 0.20705318450927734V 48080000.0ns 0.20705318450927734V 48120000.0ns 0.20705318450927734V 48600000.0ns 0.20705318450927734V 48640000.0ns 0.20705318450927734V 49360000.0ns 0.20705318450927734V 49400000.0ns 0V 49880000.0ns 0V 49920000.0ns 1.2189379930496216V 50640000.0ns 1.2189379930496216V 50680000.0ns 1.2189379930496216V 51160000.0ns 1.2189379930496216V 51200000.0ns 1.2189379930496216V 51920000.0ns 1.2189379930496216V 51960000.0ns 1.2189379930496216V 52440000.0ns 1.2189379930496216V 52480000.0ns 1.2189379930496216V 53200000.0ns 1.2189379930496216V 53240000.0ns 0V 53720000.0ns 0V 53760000.0ns 1.376880407333374V 54480000.0ns 1.376880407333374V 54520000.0ns 1.376880407333374V 55000000.0ns 1.376880407333374V 55040000.0ns 1.376880407333374V 55760000.0ns 1.376880407333374V 55800000.0ns 1.376880407333374V 56280000.0ns 1.376880407333374V 56320000.0ns 1.376880407333374V 57040000.0ns 1.376880407333374V 57080000.0ns 0V 57560000.0ns 0V 57600000.0ns 0.16451787948608398V 58320000.0ns 0.16451787948608398V 58360000.0ns 0.16451787948608398V 58840000.0ns 0.16451787948608398V 58880000.0ns 0.16451787948608398V 59600000.0ns 0.16451787948608398V 59640000.0ns 0.16451787948608398V 60120000.0ns 0.16451787948608398V 60160000.0ns 0.16451787948608398V 60880000.0ns 0.16451787948608398V 60920000.0ns 0V 61400000.0ns 0V 61440000.0ns 1.2088773250579834V 62160000.0ns 1.2088773250579834V 62200000.0ns 1.2088773250579834V 62680000.0ns 1.2088773250579834V 62720000.0ns 1.2088773250579834V 63440000.0ns 1.2088773250579834V 63480000.0ns 1.2088773250579834V 63960000.0ns 1.2088773250579834V 64000000.0ns 1.2088773250579834V 64720000.0ns 1.2088773250579834V 64760000.0ns 0V 65240000.0ns 0V 65280000.0ns 1.0731580257415771V 66000000.0ns 1.0731580257415771V 66040000.0ns 1.0731580257415771V 66520000.0ns 1.0731580257415771V 66560000.0ns 1.0731580257415771V 67280000.0ns 1.0731580257415771V 67320000.0ns 1.0731580257415771V 67800000.0ns 1.0731580257415771V 67840000.0ns 1.0731580257415771V 68560000.0ns 1.0731580257415771V 68600000.0ns 0V 69080000.0ns 0V 69120000.0ns 1.0551087856292725V 69840000.0ns 1.0551087856292725V 69880000.0ns 1.0551087856292725V 70360000.0ns 1.0551087856292725V 70400000.0ns 1.0551087856292725V 71120000.0ns 1.0551087856292725V 71160000.0ns 1.0551087856292725V 71640000.0ns 1.0551087856292725V 71680000.0ns 1.0551087856292725V 72400000.0ns 1.0551087856292725V 72440000.0ns 0V 72920000.0ns 0V 72960000.0ns 0.7520183324813843V 73680000.0ns 0.7520183324813843V 73720000.0ns 0.7520183324813843V 74200000.0ns 0.7520183324813843V 74240000.0ns 0.7520183324813843V 74960000.0ns 0.7520183324813843V 75000000.0ns 0.7520183324813843V 75480000.0ns 0.7520183324813843V 75520000.0ns 0.7520183324813843V 76240000.0ns 0.7520183324813843V 76280000.0ns 0V 76760000.0ns 0V 76800000.0ns 1.4499403238296509V 77520000.0ns 1.4499403238296509V 77560000.0ns 1.4499403238296509V 78040000.0ns 1.4499403238296509V 78080000.0ns 1.4499403238296509V 78800000.0ns 1.4499403238296509V 78840000.0ns 1.4499403238296509V 79320000.0ns 1.4499403238296509V 79360000.0ns 1.4499403238296509V 80080000.0ns 1.4499403238296509V 80120000.0ns 0V 80600000.0ns 0V 80640000.0ns 0.2956584692001343V 81360000.0ns 0.2956584692001343V 81400000.0ns 0.2956584692001343V 81880000.0ns 0.2956584692001343V 81920000.0ns 0.2956584692001343V 82640000.0ns 0.2956584692001343V 82680000.0ns 0.2956584692001343V 83160000.0ns 0.2956584692001343V 83200000.0ns 0.2956584692001343V 83920000.0ns 0.2956584692001343V 83960000.0ns 0V 84440000.0ns 0V 84480000.0ns 0.34353840351104736V 85200000.0ns 0.34353840351104736V 85240000.0ns 0.34353840351104736V 85720000.0ns 0.34353840351104736V 85760000.0ns 0.34353840351104736V 86480000.0ns 0.34353840351104736V 86520000.0ns 0.34353840351104736V 87000000.0ns 0.34353840351104736V 87040000.0ns 0.34353840351104736V 87760000.0ns 0.34353840351104736V 87800000.0ns 0V 88280000.0ns 0V 88320000.0ns 0.22561097145080566V 89040000.0ns 0.22561097145080566V 89080000.0ns 0.22561097145080566V 89560000.0ns 0.22561097145080566V 89600000.0ns 0.22561097145080566V 90320000.0ns 0.22561097145080566V 90360000.0ns 0.22561097145080566V 90840000.0ns 0.22561097145080566V 90880000.0ns 0.22561097145080566V 91600000.0ns 0.22561097145080566V 91640000.0ns 0V 92120000.0ns 0V 92160000.0ns 1.3568081855773926V 92880000.0ns 1.3568081855773926V 92920000.0ns 1.3568081855773926V 93400000.0ns 1.3568081855773926V 93440000.0ns 1.3568081855773926V 94160000.0ns 1.3568081855773926V 94200000.0ns 1.3568081855773926V 94680000.0ns 1.3568081855773926V 94720000.0ns 1.3568081855773926V 95440000.0ns 1.3568081855773926V 95480000.0ns 0V 95960000.0ns 0V 96000000.0ns 0.4793652296066284V 96720000.0ns 0.4793652296066284V 96760000.0ns 0.4793652296066284V 97240000.0ns 0.4793652296066284V 97280000.0ns 0.4793652296066284V 98000000.0ns 0.4793652296066284V 98040000.0ns 0.4793652296066284V 98520000.0ns 0.4793652296066284V 98560000.0ns 0.4793652296066284V 99280000.0ns 0.4793652296066284V 99320000.0ns 0V 99800000.0ns 0V 99840000.0ns 0.7867547273635864V 100560000.0ns 0.7867547273635864V 100600000.0ns 0.7867547273635864V 101080000.0ns 0.7867547273635864V 101120000.0ns 0.7867547273635864V 101840000.0ns 0.7867547273635864V 101880000.0ns 0.7867547273635864V 102360000.0ns 0.7867547273635864V 102400000.0ns 0.7867547273635864V 103120000.0ns 0.7867547273635864V 103160000.0ns 0V 103640000.0ns 0V 103680000.0ns 0.6138936281204224V 104400000.0ns 0.6138936281204224V 104440000.0ns 0.6138936281204224V 104920000.0ns 0.6138936281204224V 104960000.0ns 0.6138936281204224V 105680000.0ns 0.6138936281204224V 105720000.0ns 0.6138936281204224V 106200000.0ns 0.6138936281204224V 106240000.0ns 0.6138936281204224V 106960000.0ns 0.6138936281204224V 107000000.0ns 0V 107480000.0ns 0V 107520000.0ns 1.8330354690551758V 108240000.0ns 1.8330354690551758V 108280000.0ns 1.8330354690551758V 108760000.0ns 1.8330354690551758V 108800000.0ns 1.8330354690551758V 109520000.0ns 1.8330354690551758V 109560000.0ns 1.8330354690551758V 110040000.0ns 1.8330354690551758V 110080000.0ns 1.8330354690551758V 110800000.0ns 1.8330354690551758V 110840000.0ns 0V 111320000.0ns 0V 111360000.0ns 0.5352126359939575V 112080000.0ns 0.5352126359939575V 112120000.0ns 0.5352126359939575V 112600000.0ns 0.5352126359939575V 112640000.0ns 0.5352126359939575V 113360000.0ns 0.5352126359939575V 113400000.0ns 0.5352126359939575V 113880000.0ns 0.5352126359939575V 113920000.0ns 0.5352126359939575V 114640000.0ns 0.5352126359939575V 114680000.0ns 0V 115160000.0ns 0V 115200000.0ns 0.47911643981933594V 115920000.0ns 0.47911643981933594V 115960000.0ns 0.47911643981933594V 116440000.0ns 0.47911643981933594V 116480000.0ns 0.47911643981933594V 117200000.0ns 0.47911643981933594V 117240000.0ns 0.47911643981933594V 117720000.0ns 0.47911643981933594V 117760000.0ns 0.47911643981933594V 118480000.0ns 0.47911643981933594V 118520000.0ns 0V 119000000.0ns 0V 119040000.0ns 0.6288712024688721V 119760000.0ns 0.6288712024688721V 119800000.0ns 0.6288712024688721V 120280000.0ns 0.6288712024688721V 120320000.0ns 0.6288712024688721V 121040000.0ns 0.6288712024688721V 121080000.0ns 0.6288712024688721V 121560000.0ns 0.6288712024688721V 121600000.0ns 0.6288712024688721V 122320000.0ns 0.6288712024688721V 122360000.0ns 0V 122840000.0ns 0V 122880000.0ns 1.6743654012680054V 123600000.0ns 1.6743654012680054V 123640000.0ns 1.6743654012680054V 124120000.0ns 1.6743654012680054V 124160000.0ns 1.6743654012680054V 124880000.0ns 1.6743654012680054V 124920000.0ns 1.6743654012680054V 125400000.0ns 1.6743654012680054V 125440000.0ns 1.6743654012680054V 126160000.0ns 1.6743654012680054V 126200000.0ns 0V 126680000.0ns 0V 126720000.0ns 1.028953194618225V 127440000.0ns 1.028953194618225V 127480000.0ns 1.028953194618225V 127960000.0ns 1.028953194618225V 128000000.0ns 1.028953194618225V 128720000.0ns 1.028953194618225V 128760000.0ns 1.028953194618225V 129240000.0ns 1.028953194618225V 129280000.0ns 1.028953194618225V 130000000.0ns 1.028953194618225V 130040000.0ns 0V 130520000.0ns 0V 130560000.0ns 0.03515338897705078V 131280000.0ns 0.03515338897705078V 131320000.0ns 0.03515338897705078V 131800000.0ns 0.03515338897705078V 131840000.0ns 0.03515338897705078V 132560000.0ns 0.03515338897705078V 132600000.0ns 0.03515338897705078V 133080000.0ns 0.03515338897705078V 133120000.0ns 0.03515338897705078V 133840000.0ns 0.03515338897705078V 133880000.0ns 0V 134360000.0ns 0V 134400000.0ns 0.5007374286651611V 135120000.0ns 0.5007374286651611V 135160000.0ns 0.5007374286651611V 135640000.0ns 0.5007374286651611V 135680000.0ns 0.5007374286651611V 136400000.0ns 0.5007374286651611V 136440000.0ns 0.5007374286651611V 136920000.0ns 0.5007374286651611V 136960000.0ns 0.5007374286651611V 137680000.0ns 0.5007374286651611V 137720000.0ns 0V 138200000.0ns 0V 138240000.0ns 1.3598781824111938V 138960000.0ns 1.3598781824111938V 139000000.0ns 1.3598781824111938V 139480000.0ns 1.3598781824111938V 139520000.0ns 1.3598781824111938V 140240000.0ns 1.3598781824111938V 140280000.0ns 1.3598781824111938V 140760000.0ns 1.3598781824111938V 140800000.0ns 1.3598781824111938V 141520000.0ns 1.3598781824111938V 141560000.0ns 0V 142040000.0ns 0V 142080000.0ns 1.5504220724105835V 142800000.0ns 1.5504220724105835V 142840000.0ns 1.5504220724105835V 143320000.0ns 1.5504220724105835V 143360000.0ns 1.5504220724105835V 144080000.0ns 1.5504220724105835V 144120000.0ns 1.5504220724105835V 144600000.0ns 1.5504220724105835V 144640000.0ns 1.5504220724105835V 145360000.0ns 1.5504220724105835V 145400000.0ns 0V 145880000.0ns 0V 145920000.0ns 1.0550274848937988V 146640000.0ns 1.0550274848937988V 146680000.0ns 1.0550274848937988V 147160000.0ns 1.0550274848937988V 147200000.0ns 1.0550274848937988V 147920000.0ns 1.0550274848937988V 147960000.0ns 1.0550274848937988V 148440000.0ns 1.0550274848937988V 148480000.0ns 1.0550274848937988V 149200000.0ns 1.0550274848937988V 149240000.0ns 0V 149720000.0ns 0V 149760000.0ns 0.2952077388763428V 150480000.0ns 0.2952077388763428V 150520000.0ns 0.2952077388763428V 151000000.0ns 0.2952077388763428V 151040000.0ns 0.2952077388763428V 151760000.0ns 0.2952077388763428V 151800000.0ns 0.2952077388763428V 152280000.0ns 0.2952077388763428V 152320000.0ns 0.2952077388763428V 153040000.0ns 0.2952077388763428V 153080000.0ns 0V 153560000.0ns 0V 153600000.0ns 1.1526681184768677V 154320000.0ns 1.1526681184768677V 154360000.0ns 1.1526681184768677V 154840000.0ns 1.1526681184768677V 154880000.0ns 1.1526681184768677V 155600000.0ns 1.1526681184768677V 155640000.0ns 1.1526681184768677V 156120000.0ns 1.1526681184768677V 156160000.0ns 1.1526681184768677V 156880000.0ns 1.1526681184768677V 156920000.0ns 0V 157400000.0ns 0V 157440000.0ns 1.4868865013122559V 158160000.0ns 1.4868865013122559V 158200000.0ns 1.4868865013122559V 158680000.0ns 1.4868865013122559V 158720000.0ns 1.4868865013122559V 159440000.0ns 1.4868865013122559V 159480000.0ns 1.4868865013122559V 159960000.0ns 1.4868865013122559V 160000000.0ns 1.4868865013122559V 160720000.0ns 1.4868865013122559V 160760000.0ns 0V 161240000.0ns 0V 161280000.0ns 0.13019227981567383V 162000000.0ns 0.13019227981567383V 162040000.0ns 0.13019227981567383V 162520000.0ns 0.13019227981567383V 162560000.0ns 0.13019227981567383V 163280000.0ns 0.13019227981567383V 163320000.0ns 0.13019227981567383V 163800000.0ns 0.13019227981567383V 163840000.0ns 0.13019227981567383V 164560000.0ns 0.13019227981567383V 164600000.0ns 0V 165080000.0ns 0V 165120000.0ns 0.30837488174438477V 165840000.0ns 0.30837488174438477V 165880000.0ns 0.30837488174438477V 166360000.0ns 0.30837488174438477V 166400000.0ns 0.30837488174438477V 167120000.0ns 0.30837488174438477V 167160000.0ns 0.30837488174438477V 167640000.0ns 0.30837488174438477V 167680000.0ns 0.30837488174438477V 168400000.0ns 0.30837488174438477V 168440000.0ns 0V 168920000.0ns 0V 168960000.0ns 0.13420641422271729V 169680000.0ns 0.13420641422271729V 169720000.0ns 0.13420641422271729V 170200000.0ns 0.13420641422271729V 170240000.0ns 0.13420641422271729V 170960000.0ns 0.13420641422271729V 171000000.0ns 0.13420641422271729V 171480000.0ns 0.13420641422271729V 171520000.0ns 0.13420641422271729V 172240000.0ns 0.13420641422271729V 172280000.0ns 0V 172760000.0ns 0V 172800000.0ns 1.3352105617523193V 173520000.0ns 1.3352105617523193V 173560000.0ns 1.3352105617523193V 174040000.0ns 1.3352105617523193V 174080000.0ns 1.3352105617523193V 174800000.0ns 1.3352105617523193V 174840000.0ns 1.3352105617523193V 175320000.0ns 1.3352105617523193V 175360000.0ns 1.3352105617523193V 176080000.0ns 1.3352105617523193V 176120000.0ns 0V 176600000.0ns 0V 176640000.0ns 0.7921024560928345V 177360000.0ns 0.7921024560928345V 177400000.0ns 0.7921024560928345V 177880000.0ns 0.7921024560928345V 177920000.0ns 0.7921024560928345V 178640000.0ns 0.7921024560928345V 178680000.0ns 0.7921024560928345V 179160000.0ns 0.7921024560928345V 179200000.0ns 0.7921024560928345V 179920000.0ns 0.7921024560928345V 179960000.0ns 0V 180440000.0ns 0V 180480000.0ns 0.9108841419219971V 181200000.0ns 0.9108841419219971V 181240000.0ns 0.9108841419219971V 181720000.0ns 0.9108841419219971V 181760000.0ns 0.9108841419219971V 182480000.0ns 0.9108841419219971V 182520000.0ns 0.9108841419219971V 183000000.0ns 0.9108841419219971V 183040000.0ns 0.9108841419219971V 183760000.0ns 0.9108841419219971V 183800000.0ns 0V 184280000.0ns 0V 184320000.0ns 1.827146291732788V 185040000.0ns 1.827146291732788V 185080000.0ns 1.827146291732788V 185560000.0ns 1.827146291732788V 185600000.0ns 1.827146291732788V 186320000.0ns 1.827146291732788V 186360000.0ns 1.827146291732788V 186840000.0ns 1.827146291732788V 186880000.0ns 1.827146291732788V 187600000.0ns 1.827146291732788V 187640000.0ns 0V 188120000.0ns 0V 188160000.0ns 1.0180211067199707V 188880000.0ns 1.0180211067199707V 188920000.0ns 1.0180211067199707V 189400000.0ns 1.0180211067199707V 189440000.0ns 1.0180211067199707V 190160000.0ns 1.0180211067199707V 190200000.0ns 1.0180211067199707V 190680000.0ns 1.0180211067199707V 190720000.0ns 1.0180211067199707V 191440000.0ns 1.0180211067199707V 191480000.0ns 0V 191960000.0ns 0V 192000000.0ns 0.05055797100067139V 192720000.0ns 0.05055797100067139V 192760000.0ns 0.05055797100067139V 193240000.0ns 0.05055797100067139V 193280000.0ns 0.05055797100067139V 194000000.0ns 0.05055797100067139V 194040000.0ns 0.05055797100067139V 194520000.0ns 0.05055797100067139V 194560000.0ns 0.05055797100067139V 195280000.0ns 0.05055797100067139V 195320000.0ns 0V 195800000.0ns 0V 195840000.0ns 0.6037729978561401V 196560000.0ns 0.6037729978561401V 196600000.0ns 0.6037729978561401V 197080000.0ns 0.6037729978561401V 197120000.0ns 0.6037729978561401V 197840000.0ns 0.6037729978561401V 197880000.0ns 0.6037729978561401V 198360000.0ns 0.6037729978561401V 198400000.0ns 0.6037729978561401V 199120000.0ns 0.6037729978561401V 199160000.0ns 0V 199640000.0ns 0V 199680000.0ns 0.28855395317077637V 200400000.0ns 0.28855395317077637V 200440000.0ns 0.28855395317077637V 200920000.0ns 0.28855395317077637V 200960000.0ns 0.28855395317077637V 201680000.0ns 0.28855395317077637V 201720000.0ns 0.28855395317077637V 202200000.0ns 0.28855395317077637V 202240000.0ns 0.28855395317077637V 202960000.0ns 0.28855395317077637V 203000000.0ns 0V 203480000.0ns 0V 203520000.0ns 1.000589370727539V 204240000.0ns 1.000589370727539V 204280000.0ns 1.000589370727539V 204760000.0ns 1.000589370727539V 204800000.0ns 1.000589370727539V 205520000.0ns 1.000589370727539V 205560000.0ns 1.000589370727539V 206040000.0ns 1.000589370727539V 206080000.0ns 1.000589370727539V 206800000.0ns 1.000589370727539V 206840000.0ns 0V 207320000.0ns 0V 207360000.0ns 1.1583722829818726V 208080000.0ns 1.1583722829818726V 208120000.0ns 1.1583722829818726V 208600000.0ns 1.1583722829818726V 208640000.0ns 1.1583722829818726V 209360000.0ns 1.1583722829818726V 209400000.0ns 1.1583722829818726V 209880000.0ns 1.1583722829818726V 209920000.0ns 1.1583722829818726V 210640000.0ns 1.1583722829818726V 210680000.0ns 0V 211160000.0ns 0V 211200000.0ns 0.26626479625701904V 211920000.0ns 0.26626479625701904V 211960000.0ns 0.26626479625701904V 212440000.0ns 0.26626479625701904V 212480000.0ns 0.26626479625701904V 213200000.0ns 0.26626479625701904V 213240000.0ns 0.26626479625701904V 213720000.0ns 0.26626479625701904V 213760000.0ns 0.26626479625701904V 214480000.0ns 0.26626479625701904V 214520000.0ns 0V 215000000.0ns 0V 215040000.0ns 1.199228048324585V 215760000.0ns 1.199228048324585V 215800000.0ns 1.199228048324585V 216280000.0ns 1.199228048324585V 216320000.0ns 1.199228048324585V 217040000.0ns 1.199228048324585V 217080000.0ns 1.199228048324585V 217560000.0ns 1.199228048324585V 217600000.0ns 1.199228048324585V 218320000.0ns 1.199228048324585V 218360000.0ns 0V 218840000.0ns 0V 218880000.0ns 0.48730385303497314V 219600000.0ns 0.48730385303497314V 219640000.0ns 0.48730385303497314V 220120000.0ns 0.48730385303497314V 220160000.0ns 0.48730385303497314V 220880000.0ns 0.48730385303497314V 220920000.0ns 0.48730385303497314V 221400000.0ns 0.48730385303497314V 221440000.0ns 0.48730385303497314V 222160000.0ns 0.48730385303497314V 222200000.0ns 0V 222680000.0ns 0V 222720000.0ns 0.40308475494384766V 223440000.0ns 0.40308475494384766V 223480000.0ns 0.40308475494384766V 223960000.0ns 0.40308475494384766V 224000000.0ns 0.40308475494384766V 224720000.0ns 0.40308475494384766V 224760000.0ns 0.40308475494384766V 225240000.0ns 0.40308475494384766V 225280000.0ns 0.40308475494384766V 226000000.0ns 0.40308475494384766V 226040000.0ns 0V 226520000.0ns 0V 226560000.0ns 0.631257176399231V 227280000.0ns 0.631257176399231V 227320000.0ns 0.631257176399231V 227800000.0ns 0.631257176399231V 227840000.0ns 0.631257176399231V 228560000.0ns 0.631257176399231V 228600000.0ns 0.631257176399231V 229080000.0ns 0.631257176399231V 229120000.0ns 0.631257176399231V 229840000.0ns 0.631257176399231V 229880000.0ns 0V 230360000.0ns 0V 230400000.0ns 0.02771914005279541V 231120000.0ns 0.02771914005279541V 231160000.0ns 0.02771914005279541V 231640000.0ns 0.02771914005279541V 231680000.0ns 0.02771914005279541V 232400000.0ns 0.02771914005279541V 232440000.0ns 0.02771914005279541V 232920000.0ns 0.02771914005279541V 232960000.0ns 0.02771914005279541V 233680000.0ns 0.02771914005279541V 233720000.0ns 0V 234200000.0ns 0V 234240000.0ns 1.4083293676376343V 234960000.0ns 1.4083293676376343V 235000000.0ns 1.4083293676376343V 235480000.0ns 1.4083293676376343V 235520000.0ns 1.4083293676376343V 236240000.0ns 1.4083293676376343V 236280000.0ns 1.4083293676376343V 236760000.0ns 1.4083293676376343V 236800000.0ns 1.4083293676376343V 237520000.0ns 1.4083293676376343V 237560000.0ns 0V 238040000.0ns 0V 238080000.0ns 1.2673180103302002V 238800000.0ns 1.2673180103302002V 238840000.0ns 1.2673180103302002V 239320000.0ns 1.2673180103302002V 239360000.0ns 1.2673180103302002V 240080000.0ns 1.2673180103302002V 240120000.0ns 1.2673180103302002V 240600000.0ns 1.2673180103302002V 240640000.0ns 1.2673180103302002V 241360000.0ns 1.2673180103302002V 241400000.0ns 0V 241880000.0ns 0V 241920000.0ns 1.8129655122756958V 242640000.0ns 1.8129655122756958V 242680000.0ns 1.8129655122756958V 243160000.0ns 1.8129655122756958V 243200000.0ns 1.8129655122756958V 243920000.0ns 1.8129655122756958V 243960000.0ns 1.8129655122756958V 244440000.0ns 1.8129655122756958V 244480000.0ns 1.8129655122756958V 245200000.0ns 1.8129655122756958V 245240000.0ns 0V 245720000.0ns 0V 245760000.0ns 1.5064469575881958V 246480000.0ns 1.5064469575881958V 246520000.0ns 1.5064469575881958V 247000000.0ns 1.5064469575881958V 247040000.0ns 1.5064469575881958V 247760000.0ns 1.5064469575881958V 247800000.0ns 1.5064469575881958V 248280000.0ns 1.5064469575881958V 248320000.0ns 1.5064469575881958V 249040000.0ns 1.5064469575881958V 249080000.0ns 0V 249560000.0ns 0V 249600000.0ns 1.8853886127471924V 250320000.0ns 1.8853886127471924V 250360000.0ns 1.8853886127471924V 250840000.0ns 1.8853886127471924V 250880000.0ns 1.8853886127471924V 251600000.0ns 1.8853886127471924V 251640000.0ns 1.8853886127471924V 252120000.0ns 1.8853886127471924V 252160000.0ns 1.8853886127471924V 252880000.0ns 1.8853886127471924V 252920000.0ns 0V 253400000.0ns 0V 253440000.0ns 1.2043617963790894V 254160000.0ns 1.2043617963790894V 254200000.0ns 1.2043617963790894V 254680000.0ns 1.2043617963790894V 254720000.0ns 1.2043617963790894V 255440000.0ns 1.2043617963790894V 255480000.0ns 1.2043617963790894V 255960000.0ns 1.2043617963790894V 256000000.0ns 1.2043617963790894V 256720000.0ns 1.2043617963790894V 256760000.0ns 0V 257240000.0ns 0V 257280000.0ns 0.6646838188171387V 258000000.0ns 0.6646838188171387V 258040000.0ns 0.6646838188171387V 258520000.0ns 0.6646838188171387V 258560000.0ns 0.6646838188171387V 259280000.0ns 0.6646838188171387V 259320000.0ns 0.6646838188171387V 259800000.0ns 0.6646838188171387V 259840000.0ns 0.6646838188171387V 260560000.0ns 0.6646838188171387V 260600000.0ns 0V 261080000.0ns 0V 261120000.0ns 1.923681616783142V 261840000.0ns 1.923681616783142V 261880000.0ns 1.923681616783142V 262360000.0ns 1.923681616783142V 262400000.0ns 1.923681616783142V 263120000.0ns 1.923681616783142V 263160000.0ns 1.923681616783142V 263640000.0ns 1.923681616783142V 263680000.0ns 1.923681616783142V 264400000.0ns 1.923681616783142V 264440000.0ns 0V 264920000.0ns 0V 264960000.0ns 0.83675217628479V 265680000.0ns 0.83675217628479V 265720000.0ns 0.83675217628479V 266200000.0ns 0.83675217628479V 266240000.0ns 0.83675217628479V 266960000.0ns 0.83675217628479V 267000000.0ns 0.83675217628479V 267480000.0ns 0.83675217628479V 267520000.0ns 0.83675217628479V 268240000.0ns 0.83675217628479V 268280000.0ns 0V 268760000.0ns 0V 268800000.0ns 0.6513439416885376V 269520000.0ns 0.6513439416885376V 269560000.0ns 0.6513439416885376V 270040000.0ns 0.6513439416885376V 270080000.0ns 0.6513439416885376V 270800000.0ns 0.6513439416885376V 270840000.0ns 0.6513439416885376V 271320000.0ns 0.6513439416885376V 271360000.0ns 0.6513439416885376V 272080000.0ns 0.6513439416885376V 272120000.0ns 0V 272600000.0ns 0V 272640000.0ns 1.5460610389709473V 273360000.0ns 1.5460610389709473V 273400000.0ns 1.5460610389709473V 273880000.0ns 1.5460610389709473V 273920000.0ns 1.5460610389709473V 274640000.0ns 1.5460610389709473V 274680000.0ns 1.5460610389709473V 275160000.0ns 1.5460610389709473V 275200000.0ns 1.5460610389709473V 275920000.0ns 1.5460610389709473V 275960000.0ns 0V 276440000.0ns 0V 276480000.0ns 1.2786016464233398V 277200000.0ns 1.2786016464233398V 277240000.0ns 1.2786016464233398V 277720000.0ns 1.2786016464233398V 277760000.0ns 1.2786016464233398V 278480000.0ns 1.2786016464233398V 278520000.0ns 1.2786016464233398V 279000000.0ns 1.2786016464233398V 279040000.0ns 1.2786016464233398V 279760000.0ns 1.2786016464233398V 279800000.0ns 0V 280280000.0ns 0V 280320000.0ns 0.11197412014007568V 281040000.0ns 0.11197412014007568V 281080000.0ns 0.11197412014007568V 281560000.0ns 0.11197412014007568V 281600000.0ns 0.11197412014007568V 282320000.0ns 0.11197412014007568V 282360000.0ns 0.11197412014007568V 282840000.0ns 0.11197412014007568V 282880000.0ns 0.11197412014007568V 283600000.0ns 0.11197412014007568V 283640000.0ns 0V 284120000.0ns 0V 284160000.0ns 1.5291328430175781V 284880000.0ns 1.5291328430175781V 284920000.0ns 1.5291328430175781V 285400000.0ns 1.5291328430175781V 285440000.0ns 1.5291328430175781V 286160000.0ns 1.5291328430175781V 286200000.0ns 1.5291328430175781V 286680000.0ns 1.5291328430175781V 286720000.0ns 1.5291328430175781V 287440000.0ns 1.5291328430175781V 287480000.0ns 0V 287960000.0ns 0V 288000000.0ns 1.028652310371399V 288720000.0ns 1.028652310371399V 288760000.0ns 1.028652310371399V 289240000.0ns 1.028652310371399V 289280000.0ns 1.028652310371399V 290000000.0ns 1.028652310371399V 290040000.0ns 1.028652310371399V 290520000.0ns 1.028652310371399V 290560000.0ns 1.028652310371399V 291280000.0ns 1.028652310371399V 291320000.0ns 0V 291800000.0ns 0V 291840000.0ns 0.9055479764938354V 292560000.0ns 0.9055479764938354V 292600000.0ns 0.9055479764938354V 293080000.0ns 0.9055479764938354V 293120000.0ns 0.9055479764938354V 293840000.0ns 0.9055479764938354V 293880000.0ns 0.9055479764938354V 294360000.0ns 0.9055479764938354V 294400000.0ns 0.9055479764938354V 295120000.0ns 0.9055479764938354V 295160000.0ns 0V 295640000.0ns 0V 295680000.0ns 0.7932971715927124V 296400000.0ns 0.7932971715927124V 296440000.0ns 0.7932971715927124V 296920000.0ns 0.7932971715927124V 296960000.0ns 0.7932971715927124V 297680000.0ns 0.7932971715927124V 297720000.0ns 0.7932971715927124V 298200000.0ns 0.7932971715927124V 298240000.0ns 0.7932971715927124V 298960000.0ns 0.7932971715927124V 299000000.0ns 0V 299480000.0ns 0V 299520000.0ns 0.021576762199401855V 300240000.0ns 0.021576762199401855V 300280000.0ns 0.021576762199401855V 300760000.0ns 0.021576762199401855V 300800000.0ns 0.021576762199401855V 301520000.0ns 0.021576762199401855V 301560000.0ns 0.021576762199401855V 302040000.0ns 0.021576762199401855V 302080000.0ns 0.021576762199401855V 302800000.0ns 0.021576762199401855V 302840000.0ns 0V 303320000.0ns 0V 303360000.0ns 1.1066228151321411V 304080000.0ns 1.1066228151321411V 304120000.0ns 1.1066228151321411V 304600000.0ns 1.1066228151321411V 304640000.0ns 1.1066228151321411V 305360000.0ns 1.1066228151321411V 305400000.0ns 1.1066228151321411V 305880000.0ns 1.1066228151321411V 305920000.0ns 1.1066228151321411V 306640000.0ns 1.1066228151321411V 306680000.0ns 0V 307160000.0ns 0V 307200000.0ns 0.41128110885620117V 307920000.0ns 0.41128110885620117V 307960000.0ns 0.41128110885620117V 308440000.0ns 0.41128110885620117V 308480000.0ns 0.41128110885620117V 309200000.0ns 0.41128110885620117V 309240000.0ns 0.41128110885620117V 309720000.0ns 0.41128110885620117V 309760000.0ns 0.41128110885620117V 310480000.0ns 0.41128110885620117V 310520000.0ns 0V 311000000.0ns 0V 311040000.0ns 0.411934494972229V 311760000.0ns 0.411934494972229V 311800000.0ns 0.411934494972229V 312280000.0ns 0.411934494972229V 312320000.0ns 0.411934494972229V 313040000.0ns 0.411934494972229V 313080000.0ns 0.411934494972229V 313560000.0ns 0.411934494972229V 313600000.0ns 0.411934494972229V 314320000.0ns 0.411934494972229V 314360000.0ns 0V 314840000.0ns 0V 314880000.0ns 0.8076795339584351V 315600000.0ns 0.8076795339584351V 315640000.0ns 0.8076795339584351V 316120000.0ns 0.8076795339584351V 316160000.0ns 0.8076795339584351V 316880000.0ns 0.8076795339584351V 316920000.0ns 0.8076795339584351V 317400000.0ns 0.8076795339584351V 317440000.0ns 0.8076795339584351V 318160000.0ns 0.8076795339584351V 318200000.0ns 0V 318680000.0ns 0V 318720000.0ns 1.239526391029358V 319440000.0ns 1.239526391029358V 319480000.0ns 1.239526391029358V 319960000.0ns 1.239526391029358V 320000000.0ns 1.239526391029358V 320720000.0ns 1.239526391029358V 320760000.0ns 1.239526391029358V 321240000.0ns 1.239526391029358V 321280000.0ns 1.239526391029358V 322000000.0ns 1.239526391029358V 322040000.0ns 0V 322520000.0ns 0V 322560000.0ns 0.8498064279556274V 323280000.0ns 0.8498064279556274V 323320000.0ns 0.8498064279556274V 323800000.0ns 0.8498064279556274V 323840000.0ns 0.8498064279556274V 324560000.0ns 0.8498064279556274V 324600000.0ns 0.8498064279556274V 325080000.0ns 0.8498064279556274V 325120000.0ns 0.8498064279556274V 325840000.0ns 0.8498064279556274V 325880000.0ns 0V 326360000.0ns 0V 326400000.0ns 1.2954885959625244V 327120000.0ns 1.2954885959625244V 327160000.0ns 1.2954885959625244V 327640000.0ns 1.2954885959625244V 327680000.0ns 1.2954885959625244V 328400000.0ns 1.2954885959625244V 328440000.0ns 1.2954885959625244V 328920000.0ns 1.2954885959625244V 328960000.0ns 1.2954885959625244V 329680000.0ns 1.2954885959625244V 329720000.0ns 0V 330200000.0ns 0V 330240000.0ns 1.5997889041900635V 330960000.0ns 1.5997889041900635V 331000000.0ns 1.5997889041900635V 331480000.0ns 1.5997889041900635V 331520000.0ns 1.5997889041900635V 332240000.0ns 1.5997889041900635V 332280000.0ns 1.5997889041900635V 332760000.0ns 1.5997889041900635V 332800000.0ns 1.5997889041900635V 333520000.0ns 1.5997889041900635V 333560000.0ns 0V 334040000.0ns 0V 334080000.0ns 0.7632800340652466V 334800000.0ns 0.7632800340652466V 334840000.0ns 0.7632800340652466V 335320000.0ns 0.7632800340652466V 335360000.0ns 0.7632800340652466V 336080000.0ns 0.7632800340652466V 336120000.0ns 0.7632800340652466V 336600000.0ns 0.7632800340652466V 336640000.0ns 0.7632800340652466V 337360000.0ns 0.7632800340652466V 337400000.0ns 0V 337880000.0ns 0V 337920000.0ns 0.05809962749481201V 338640000.0ns 0.05809962749481201V 338680000.0ns 0.05809962749481201V 339160000.0ns 0.05809962749481201V 339200000.0ns 0.05809962749481201V 339920000.0ns 0.05809962749481201V 339960000.0ns 0.05809962749481201V 340440000.0ns 0.05809962749481201V 340480000.0ns 0.05809962749481201V 341200000.0ns 0.05809962749481201V 341240000.0ns 0V 341720000.0ns 0V 341760000.0ns 1.4315754175186157V 342480000.0ns 1.4315754175186157V 342520000.0ns 1.4315754175186157V 343000000.0ns 1.4315754175186157V 343040000.0ns 1.4315754175186157V 343760000.0ns 1.4315754175186157V 343800000.0ns 1.4315754175186157V 344280000.0ns 1.4315754175186157V 344320000.0ns 1.4315754175186157V 345040000.0ns 1.4315754175186157V 345080000.0ns 0V 345560000.0ns 0V 345600000.0ns 1.662571907043457V 346320000.0ns 1.662571907043457V 346360000.0ns 1.662571907043457V 346840000.0ns 1.662571907043457V 346880000.0ns 1.662571907043457V 347600000.0ns 1.662571907043457V 347640000.0ns 1.662571907043457V 348120000.0ns 1.662571907043457V 348160000.0ns 1.662571907043457V 348880000.0ns 1.662571907043457V 348920000.0ns 0V 349400000.0ns 0V 349440000.0ns 0.8203641176223755V 350160000.0ns 0.8203641176223755V 350200000.0ns 0.8203641176223755V 350680000.0ns 0.8203641176223755V 350720000.0ns 0.8203641176223755V 351440000.0ns 0.8203641176223755V 351480000.0ns 0.8203641176223755V 351960000.0ns 0.8203641176223755V 352000000.0ns 0.8203641176223755V 352720000.0ns 0.8203641176223755V 352760000.0ns 0V 353240000.0ns 0V 353280000.0ns 1.6321138143539429V 354000000.0ns 1.6321138143539429V 354040000.0ns 1.6321138143539429V 354520000.0ns 1.6321138143539429V 354560000.0ns 1.6321138143539429V 355280000.0ns 1.6321138143539429V 355320000.0ns 1.6321138143539429V 355800000.0ns 1.6321138143539429V 355840000.0ns 1.6321138143539429V 356560000.0ns 1.6321138143539429V 356600000.0ns 0V 357080000.0ns 0V 357120000.0ns 0.5078330039978027V 357840000.0ns 0.5078330039978027V 357880000.0ns 0.5078330039978027V 358360000.0ns 0.5078330039978027V 358400000.0ns 0.5078330039978027V 359120000.0ns 0.5078330039978027V 359160000.0ns 0.5078330039978027V 359640000.0ns 0.5078330039978027V 359680000.0ns 0.5078330039978027V 360400000.0ns 0.5078330039978027V 360440000.0ns 0V 360920000.0ns 0V 360960000.0ns 0.5386412143707275V 361680000.0ns 0.5386412143707275V 361720000.0ns 0.5386412143707275V 362200000.0ns 0.5386412143707275V 362240000.0ns 0.5386412143707275V 362960000.0ns 0.5386412143707275V 363000000.0ns 0.5386412143707275V 363480000.0ns 0.5386412143707275V 363520000.0ns 0.5386412143707275V 364240000.0ns 0.5386412143707275V 364280000.0ns 0V 364760000.0ns 0V 364800000.0ns 0.9434295892715454V 365520000.0ns 0.9434295892715454V 365560000.0ns 0.9434295892715454V 366040000.0ns 0.9434295892715454V 366080000.0ns 0.9434295892715454V 366800000.0ns 0.9434295892715454V 366840000.0ns 0.9434295892715454V 367320000.0ns 0.9434295892715454V 367360000.0ns 0.9434295892715454V 368080000.0ns 0.9434295892715454V 368120000.0ns 0V 368600000.0ns 0V 368640000.0ns 1.6125825643539429V 369360000.0ns 1.6125825643539429V 369400000.0ns 1.6125825643539429V 369880000.0ns 1.6125825643539429V 369920000.0ns 1.6125825643539429V 370640000.0ns 1.6125825643539429V 370680000.0ns 1.6125825643539429V 371160000.0ns 1.6125825643539429V 371200000.0ns 1.6125825643539429V 371920000.0ns 1.6125825643539429V 371960000.0ns 0V 372440000.0ns 0V 372480000.0ns 1.1577459573745728V 373200000.0ns 1.1577459573745728V 373240000.0ns 1.1577459573745728V 373720000.0ns 1.1577459573745728V 373760000.0ns 1.1577459573745728V 374480000.0ns 1.1577459573745728V 374520000.0ns 1.1577459573745728V 375000000.0ns 1.1577459573745728V 375040000.0ns 1.1577459573745728V 375760000.0ns 1.1577459573745728V 375800000.0ns 0V 376280000.0ns 0V 376320000.0ns 1.9656106233596802V 377040000.0ns 1.9656106233596802V 377080000.0ns 1.9656106233596802V 377560000.0ns 1.9656106233596802V 377600000.0ns 1.9656106233596802V 378320000.0ns 1.9656106233596802V 378360000.0ns 1.9656106233596802V 378840000.0ns 1.9656106233596802V 378880000.0ns 1.9656106233596802V 379600000.0ns 1.9656106233596802V 379640000.0ns 0V 380120000.0ns 0V 380160000.0ns 1.1139044761657715V 380880000.0ns 1.1139044761657715V 380920000.0ns 1.1139044761657715V 381400000.0ns 1.1139044761657715V 381440000.0ns 1.1139044761657715V 382160000.0ns 1.1139044761657715V 382200000.0ns 1.1139044761657715V 382680000.0ns 1.1139044761657715V 382720000.0ns 1.1139044761657715V 383440000.0ns 1.1139044761657715V 383480000.0ns 0V 383960000.0ns 0V 384000000.0ns 1.2732863426208496V 384720000.0ns 1.2732863426208496V 384760000.0ns 1.2732863426208496V 385240000.0ns 1.2732863426208496V 385280000.0ns 1.2732863426208496V 386000000.0ns 1.2732863426208496V 386040000.0ns 1.2732863426208496V 386520000.0ns 1.2732863426208496V 386560000.0ns 1.2732863426208496V 387280000.0ns 1.2732863426208496V 387320000.0ns 0V 387800000.0ns 0V 387840000.0ns 1.6230039596557617V 388560000.0ns 1.6230039596557617V 388600000.0ns 1.6230039596557617V 389080000.0ns 1.6230039596557617V 389120000.0ns 1.6230039596557617V 389840000.0ns 1.6230039596557617V 389880000.0ns 1.6230039596557617V 390360000.0ns 1.6230039596557617V 390400000.0ns 1.6230039596557617V 391120000.0ns 1.6230039596557617V 391160000.0ns 0V)
VX_1 X_1 0 PWL(0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 1.8190712928771973V 8400000.0ns 1.8190712928771973V 8440000.0ns 1.8190712928771973V 8920000.0ns 1.8190712928771973V 8960000.0ns 1.8190712928771973V 9680000.0ns 1.8190712928771973V 9720000.0ns 1.8190712928771973V 10200000.0ns 1.8190712928771973V 10240000.0ns 1.8190712928771973V 10960000.0ns 1.8190712928771973V 11000000.0ns 0V 11480000.0ns 0V 11520000.0ns 1.6753596067428589V 12240000.0ns 1.6753596067428589V 12280000.0ns 1.6753596067428589V 12760000.0ns 1.6753596067428589V 12800000.0ns 1.6753596067428589V 13520000.0ns 1.6753596067428589V 13560000.0ns 1.6753596067428589V 14040000.0ns 1.6753596067428589V 14080000.0ns 1.6753596067428589V 14800000.0ns 1.6753596067428589V 14840000.0ns 0V 15320000.0ns 0V 15360000.0ns 0.027140378952026367V 16080000.0ns 0.027140378952026367V 16120000.0ns 0.027140378952026367V 16600000.0ns 0.027140378952026367V 16640000.0ns 0.027140378952026367V 17360000.0ns 0.027140378952026367V 17400000.0ns 0.027140378952026367V 17880000.0ns 0.027140378952026367V 17920000.0ns 0.027140378952026367V 18640000.0ns 0.027140378952026367V 18680000.0ns 0V 19160000.0ns 0V 19200000.0ns 1.0674731731414795V 19920000.0ns 1.0674731731414795V 19960000.0ns 1.0674731731414795V 20440000.0ns 1.0674731731414795V 20480000.0ns 1.0674731731414795V 21200000.0ns 1.0674731731414795V 21240000.0ns 1.0674731731414795V 21720000.0ns 1.0674731731414795V 21760000.0ns 1.0674731731414795V 22480000.0ns 1.0674731731414795V 22520000.0ns 0V 23000000.0ns 0V 23040000.0ns 1.611703872680664V 23760000.0ns 1.611703872680664V 23800000.0ns 1.611703872680664V 24280000.0ns 1.611703872680664V 24320000.0ns 1.611703872680664V 25040000.0ns 1.611703872680664V 25080000.0ns 1.611703872680664V 25560000.0ns 1.611703872680664V 25600000.0ns 1.611703872680664V 26320000.0ns 1.611703872680664V 26360000.0ns 0V 26840000.0ns 0V 26880000.0ns 0.1788259744644165V 27600000.0ns 0.1788259744644165V 27640000.0ns 0.1788259744644165V 28120000.0ns 0.1788259744644165V 28160000.0ns 0.1788259744644165V 28880000.0ns 0.1788259744644165V 28920000.0ns 0.1788259744644165V 29400000.0ns 0.1788259744644165V 29440000.0ns 0.1788259744644165V 30160000.0ns 0.1788259744644165V 30200000.0ns 0V 30680000.0ns 0V 30720000.0ns 0.6219770908355713V 31440000.0ns 0.6219770908355713V 31480000.0ns 0.6219770908355713V 31960000.0ns 0.6219770908355713V 32000000.0ns 0.6219770908355713V 32720000.0ns 0.6219770908355713V 32760000.0ns 0.6219770908355713V 33240000.0ns 0.6219770908355713V 33280000.0ns 0.6219770908355713V 34000000.0ns 0.6219770908355713V 34040000.0ns 0V 34520000.0ns 0V 34560000.0ns 0.026337623596191406V 35280000.0ns 0.026337623596191406V 35320000.0ns 0.026337623596191406V 35800000.0ns 0.026337623596191406V 35840000.0ns 0.026337623596191406V 36560000.0ns 0.026337623596191406V 36600000.0ns 0.026337623596191406V 37080000.0ns 0.026337623596191406V 37120000.0ns 0.026337623596191406V 37840000.0ns 0.026337623596191406V 37880000.0ns 0V 38360000.0ns 0V 38400000.0ns 1.9300395250320435V 39120000.0ns 1.9300395250320435V 39160000.0ns 1.9300395250320435V 39640000.0ns 1.9300395250320435V 39680000.0ns 1.9300395250320435V 40400000.0ns 1.9300395250320435V 40440000.0ns 1.9300395250320435V 40920000.0ns 1.9300395250320435V 40960000.0ns 1.9300395250320435V 41680000.0ns 1.9300395250320435V 41720000.0ns 0V 42200000.0ns 0V 42240000.0ns 1.5200536251068115V 42960000.0ns 1.5200536251068115V 43000000.0ns 1.5200536251068115V 43480000.0ns 1.5200536251068115V 43520000.0ns 1.5200536251068115V 44240000.0ns 1.5200536251068115V 44280000.0ns 1.5200536251068115V 44760000.0ns 1.5200536251068115V 44800000.0ns 1.5200536251068115V 45520000.0ns 1.5200536251068115V 45560000.0ns 0V 46040000.0ns 0V 46080000.0ns 1.7929468154907227V 46800000.0ns 1.7929468154907227V 46840000.0ns 1.7929468154907227V 47320000.0ns 1.7929468154907227V 47360000.0ns 1.7929468154907227V 48080000.0ns 1.7929468154907227V 48120000.0ns 1.7929468154907227V 48600000.0ns 1.7929468154907227V 48640000.0ns 1.7929468154907227V 49360000.0ns 1.7929468154907227V 49400000.0ns 0V 49880000.0ns 0V 49920000.0ns 0.7810620069503784V 50640000.0ns 0.7810620069503784V 50680000.0ns 0.7810620069503784V 51160000.0ns 0.7810620069503784V 51200000.0ns 0.7810620069503784V 51920000.0ns 0.7810620069503784V 51960000.0ns 0.7810620069503784V 52440000.0ns 0.7810620069503784V 52480000.0ns 0.7810620069503784V 53200000.0ns 0.7810620069503784V 53240000.0ns 0V 53720000.0ns 0V 53760000.0ns 0.623119592666626V 54480000.0ns 0.623119592666626V 54520000.0ns 0.623119592666626V 55000000.0ns 0.623119592666626V 55040000.0ns 0.623119592666626V 55760000.0ns 0.623119592666626V 55800000.0ns 0.623119592666626V 56280000.0ns 0.623119592666626V 56320000.0ns 0.623119592666626V 57040000.0ns 0.623119592666626V 57080000.0ns 0V 57560000.0ns 0V 57600000.0ns 1.835482120513916V 58320000.0ns 1.835482120513916V 58360000.0ns 1.835482120513916V 58840000.0ns 1.835482120513916V 58880000.0ns 1.835482120513916V 59600000.0ns 1.835482120513916V 59640000.0ns 1.835482120513916V 60120000.0ns 1.835482120513916V 60160000.0ns 1.835482120513916V 60880000.0ns 1.835482120513916V 60920000.0ns 0V 61400000.0ns 0V 61440000.0ns 0.7911226749420166V 62160000.0ns 0.7911226749420166V 62200000.0ns 0.7911226749420166V 62680000.0ns 0.7911226749420166V 62720000.0ns 0.7911226749420166V 63440000.0ns 0.7911226749420166V 63480000.0ns 0.7911226749420166V 63960000.0ns 0.7911226749420166V 64000000.0ns 0.7911226749420166V 64720000.0ns 0.7911226749420166V 64760000.0ns 0V 65240000.0ns 0V 65280000.0ns 0.9268419742584229V 66000000.0ns 0.9268419742584229V 66040000.0ns 0.9268419742584229V 66520000.0ns 0.9268419742584229V 66560000.0ns 0.9268419742584229V 67280000.0ns 0.9268419742584229V 67320000.0ns 0.9268419742584229V 67800000.0ns 0.9268419742584229V 67840000.0ns 0.9268419742584229V 68560000.0ns 0.9268419742584229V 68600000.0ns 0V 69080000.0ns 0V 69120000.0ns 0.9448912143707275V 69840000.0ns 0.9448912143707275V 69880000.0ns 0.9448912143707275V 70360000.0ns 0.9448912143707275V 70400000.0ns 0.9448912143707275V 71120000.0ns 0.9448912143707275V 71160000.0ns 0.9448912143707275V 71640000.0ns 0.9448912143707275V 71680000.0ns 0.9448912143707275V 72400000.0ns 0.9448912143707275V 72440000.0ns 0V 72920000.0ns 0V 72960000.0ns 1.2479816675186157V 73680000.0ns 1.2479816675186157V 73720000.0ns 1.2479816675186157V 74200000.0ns 1.2479816675186157V 74240000.0ns 1.2479816675186157V 74960000.0ns 1.2479816675186157V 75000000.0ns 1.2479816675186157V 75480000.0ns 1.2479816675186157V 75520000.0ns 1.2479816675186157V 76240000.0ns 1.2479816675186157V 76280000.0ns 0V 76760000.0ns 0V 76800000.0ns 0.5500596761703491V 77520000.0ns 0.5500596761703491V 77560000.0ns 0.5500596761703491V 78040000.0ns 0.5500596761703491V 78080000.0ns 0.5500596761703491V 78800000.0ns 0.5500596761703491V 78840000.0ns 0.5500596761703491V 79320000.0ns 0.5500596761703491V 79360000.0ns 0.5500596761703491V 80080000.0ns 0.5500596761703491V 80120000.0ns 0V 80600000.0ns 0V 80640000.0ns 1.7043415307998657V 81360000.0ns 1.7043415307998657V 81400000.0ns 1.7043415307998657V 81880000.0ns 1.7043415307998657V 81920000.0ns 1.7043415307998657V 82640000.0ns 1.7043415307998657V 82680000.0ns 1.7043415307998657V 83160000.0ns 1.7043415307998657V 83200000.0ns 1.7043415307998657V 83920000.0ns 1.7043415307998657V 83960000.0ns 0V 84440000.0ns 0V 84480000.0ns 1.6564615964889526V 85200000.0ns 1.6564615964889526V 85240000.0ns 1.6564615964889526V 85720000.0ns 1.6564615964889526V 85760000.0ns 1.6564615964889526V 86480000.0ns 1.6564615964889526V 86520000.0ns 1.6564615964889526V 87000000.0ns 1.6564615964889526V 87040000.0ns 1.6564615964889526V 87760000.0ns 1.6564615964889526V 87800000.0ns 0V 88280000.0ns 0V 88320000.0ns 1.7743890285491943V 89040000.0ns 1.7743890285491943V 89080000.0ns 1.7743890285491943V 89560000.0ns 1.7743890285491943V 89600000.0ns 1.7743890285491943V 90320000.0ns 1.7743890285491943V 90360000.0ns 1.7743890285491943V 90840000.0ns 1.7743890285491943V 90880000.0ns 1.7743890285491943V 91600000.0ns 1.7743890285491943V 91640000.0ns 0V 92120000.0ns 0V 92160000.0ns 0.6431918144226074V 92880000.0ns 0.6431918144226074V 92920000.0ns 0.6431918144226074V 93400000.0ns 0.6431918144226074V 93440000.0ns 0.6431918144226074V 94160000.0ns 0.6431918144226074V 94200000.0ns 0.6431918144226074V 94680000.0ns 0.6431918144226074V 94720000.0ns 0.6431918144226074V 95440000.0ns 0.6431918144226074V 95480000.0ns 0V 95960000.0ns 0V 96000000.0ns 1.5206347703933716V 96720000.0ns 1.5206347703933716V 96760000.0ns 1.5206347703933716V 97240000.0ns 1.5206347703933716V 97280000.0ns 1.5206347703933716V 98000000.0ns 1.5206347703933716V 98040000.0ns 1.5206347703933716V 98520000.0ns 1.5206347703933716V 98560000.0ns 1.5206347703933716V 99280000.0ns 1.5206347703933716V 99320000.0ns 0V 99800000.0ns 0V 99840000.0ns 1.2132452726364136V 100560000.0ns 1.2132452726364136V 100600000.0ns 1.2132452726364136V 101080000.0ns 1.2132452726364136V 101120000.0ns 1.2132452726364136V 101840000.0ns 1.2132452726364136V 101880000.0ns 1.2132452726364136V 102360000.0ns 1.2132452726364136V 102400000.0ns 1.2132452726364136V 103120000.0ns 1.2132452726364136V 103160000.0ns 0V 103640000.0ns 0V 103680000.0ns 1.3861063718795776V 104400000.0ns 1.3861063718795776V 104440000.0ns 1.3861063718795776V 104920000.0ns 1.3861063718795776V 104960000.0ns 1.3861063718795776V 105680000.0ns 1.3861063718795776V 105720000.0ns 1.3861063718795776V 106200000.0ns 1.3861063718795776V 106240000.0ns 1.3861063718795776V 106960000.0ns 1.3861063718795776V 107000000.0ns 0V 107480000.0ns 0V 107520000.0ns 0.16696453094482422V 108240000.0ns 0.16696453094482422V 108280000.0ns 0.16696453094482422V 108760000.0ns 0.16696453094482422V 108800000.0ns 0.16696453094482422V 109520000.0ns 0.16696453094482422V 109560000.0ns 0.16696453094482422V 110040000.0ns 0.16696453094482422V 110080000.0ns 0.16696453094482422V 110800000.0ns 0.16696453094482422V 110840000.0ns 0V 111320000.0ns 0V 111360000.0ns 1.4647873640060425V 112080000.0ns 1.4647873640060425V 112120000.0ns 1.4647873640060425V 112600000.0ns 1.4647873640060425V 112640000.0ns 1.4647873640060425V 113360000.0ns 1.4647873640060425V 113400000.0ns 1.4647873640060425V 113880000.0ns 1.4647873640060425V 113920000.0ns 1.4647873640060425V 114640000.0ns 1.4647873640060425V 114680000.0ns 0V 115160000.0ns 0V 115200000.0ns 1.520883560180664V 115920000.0ns 1.520883560180664V 115960000.0ns 1.520883560180664V 116440000.0ns 1.520883560180664V 116480000.0ns 1.520883560180664V 117200000.0ns 1.520883560180664V 117240000.0ns 1.520883560180664V 117720000.0ns 1.520883560180664V 117760000.0ns 1.520883560180664V 118480000.0ns 1.520883560180664V 118520000.0ns 0V 119000000.0ns 0V 119040000.0ns 1.371128797531128V 119760000.0ns 1.371128797531128V 119800000.0ns 1.371128797531128V 120280000.0ns 1.371128797531128V 120320000.0ns 1.371128797531128V 121040000.0ns 1.371128797531128V 121080000.0ns 1.371128797531128V 121560000.0ns 1.371128797531128V 121600000.0ns 1.371128797531128V 122320000.0ns 1.371128797531128V 122360000.0ns 0V 122840000.0ns 0V 122880000.0ns 0.32563459873199463V 123600000.0ns 0.32563459873199463V 123640000.0ns 0.32563459873199463V 124120000.0ns 0.32563459873199463V 124160000.0ns 0.32563459873199463V 124880000.0ns 0.32563459873199463V 124920000.0ns 0.32563459873199463V 125400000.0ns 0.32563459873199463V 125440000.0ns 0.32563459873199463V 126160000.0ns 0.32563459873199463V 126200000.0ns 0V 126680000.0ns 0V 126720000.0ns 0.9710468053817749V 127440000.0ns 0.9710468053817749V 127480000.0ns 0.9710468053817749V 127960000.0ns 0.9710468053817749V 128000000.0ns 0.9710468053817749V 128720000.0ns 0.9710468053817749V 128760000.0ns 0.9710468053817749V 129240000.0ns 0.9710468053817749V 129280000.0ns 0.9710468053817749V 130000000.0ns 0.9710468053817749V 130040000.0ns 0V 130520000.0ns 0V 130560000.0ns 1.9648466110229492V 131280000.0ns 1.9648466110229492V 131320000.0ns 1.9648466110229492V 131800000.0ns 1.9648466110229492V 131840000.0ns 1.9648466110229492V 132560000.0ns 1.9648466110229492V 132600000.0ns 1.9648466110229492V 133080000.0ns 1.9648466110229492V 133120000.0ns 1.9648466110229492V 133840000.0ns 1.9648466110229492V 133880000.0ns 0V 134360000.0ns 0V 134400000.0ns 1.4992625713348389V 135120000.0ns 1.4992625713348389V 135160000.0ns 1.4992625713348389V 135640000.0ns 1.4992625713348389V 135680000.0ns 1.4992625713348389V 136400000.0ns 1.4992625713348389V 136440000.0ns 1.4992625713348389V 136920000.0ns 1.4992625713348389V 136960000.0ns 1.4992625713348389V 137680000.0ns 1.4992625713348389V 137720000.0ns 0V 138200000.0ns 0V 138240000.0ns 0.6401218175888062V 138960000.0ns 0.6401218175888062V 139000000.0ns 0.6401218175888062V 139480000.0ns 0.6401218175888062V 139520000.0ns 0.6401218175888062V 140240000.0ns 0.6401218175888062V 140280000.0ns 0.6401218175888062V 140760000.0ns 0.6401218175888062V 140800000.0ns 0.6401218175888062V 141520000.0ns 0.6401218175888062V 141560000.0ns 0V 142040000.0ns 0V 142080000.0ns 0.4495779275894165V 142800000.0ns 0.4495779275894165V 142840000.0ns 0.4495779275894165V 143320000.0ns 0.4495779275894165V 143360000.0ns 0.4495779275894165V 144080000.0ns 0.4495779275894165V 144120000.0ns 0.4495779275894165V 144600000.0ns 0.4495779275894165V 144640000.0ns 0.4495779275894165V 145360000.0ns 0.4495779275894165V 145400000.0ns 0V 145880000.0ns 0V 145920000.0ns 0.9449725151062012V 146640000.0ns 0.9449725151062012V 146680000.0ns 0.9449725151062012V 147160000.0ns 0.9449725151062012V 147200000.0ns 0.9449725151062012V 147920000.0ns 0.9449725151062012V 147960000.0ns 0.9449725151062012V 148440000.0ns 0.9449725151062012V 148480000.0ns 0.9449725151062012V 149200000.0ns 0.9449725151062012V 149240000.0ns 0V 149720000.0ns 0V 149760000.0ns 1.7047922611236572V 150480000.0ns 1.7047922611236572V 150520000.0ns 1.7047922611236572V 151000000.0ns 1.7047922611236572V 151040000.0ns 1.7047922611236572V 151760000.0ns 1.7047922611236572V 151800000.0ns 1.7047922611236572V 152280000.0ns 1.7047922611236572V 152320000.0ns 1.7047922611236572V 153040000.0ns 1.7047922611236572V 153080000.0ns 0V 153560000.0ns 0V 153600000.0ns 0.8473318815231323V 154320000.0ns 0.8473318815231323V 154360000.0ns 0.8473318815231323V 154840000.0ns 0.8473318815231323V 154880000.0ns 0.8473318815231323V 155600000.0ns 0.8473318815231323V 155640000.0ns 0.8473318815231323V 156120000.0ns 0.8473318815231323V 156160000.0ns 0.8473318815231323V 156880000.0ns 0.8473318815231323V 156920000.0ns 0V 157400000.0ns 0V 157440000.0ns 0.5131134986877441V 158160000.0ns 0.5131134986877441V 158200000.0ns 0.5131134986877441V 158680000.0ns 0.5131134986877441V 158720000.0ns 0.5131134986877441V 159440000.0ns 0.5131134986877441V 159480000.0ns 0.5131134986877441V 159960000.0ns 0.5131134986877441V 160000000.0ns 0.5131134986877441V 160720000.0ns 0.5131134986877441V 160760000.0ns 0V 161240000.0ns 0V 161280000.0ns 1.8698077201843262V 162000000.0ns 1.8698077201843262V 162040000.0ns 1.8698077201843262V 162520000.0ns 1.8698077201843262V 162560000.0ns 1.8698077201843262V 163280000.0ns 1.8698077201843262V 163320000.0ns 1.8698077201843262V 163800000.0ns 1.8698077201843262V 163840000.0ns 1.8698077201843262V 164560000.0ns 1.8698077201843262V 164600000.0ns 0V 165080000.0ns 0V 165120000.0ns 1.6916251182556152V 165840000.0ns 1.6916251182556152V 165880000.0ns 1.6916251182556152V 166360000.0ns 1.6916251182556152V 166400000.0ns 1.6916251182556152V 167120000.0ns 1.6916251182556152V 167160000.0ns 1.6916251182556152V 167640000.0ns 1.6916251182556152V 167680000.0ns 1.6916251182556152V 168400000.0ns 1.6916251182556152V 168440000.0ns 0V 168920000.0ns 0V 168960000.0ns 1.8657935857772827V 169680000.0ns 1.8657935857772827V 169720000.0ns 1.8657935857772827V 170200000.0ns 1.8657935857772827V 170240000.0ns 1.8657935857772827V 170960000.0ns 1.8657935857772827V 171000000.0ns 1.8657935857772827V 171480000.0ns 1.8657935857772827V 171520000.0ns 1.8657935857772827V 172240000.0ns 1.8657935857772827V 172280000.0ns 0V 172760000.0ns 0V 172800000.0ns 0.6647894382476807V 173520000.0ns 0.6647894382476807V 173560000.0ns 0.6647894382476807V 174040000.0ns 0.6647894382476807V 174080000.0ns 0.6647894382476807V 174800000.0ns 0.6647894382476807V 174840000.0ns 0.6647894382476807V 175320000.0ns 0.6647894382476807V 175360000.0ns 0.6647894382476807V 176080000.0ns 0.6647894382476807V 176120000.0ns 0V 176600000.0ns 0V 176640000.0ns 1.2078975439071655V 177360000.0ns 1.2078975439071655V 177400000.0ns 1.2078975439071655V 177880000.0ns 1.2078975439071655V 177920000.0ns 1.2078975439071655V 178640000.0ns 1.2078975439071655V 178680000.0ns 1.2078975439071655V 179160000.0ns 1.2078975439071655V 179200000.0ns 1.2078975439071655V 179920000.0ns 1.2078975439071655V 179960000.0ns 0V 180440000.0ns 0V 180480000.0ns 1.089115858078003V 181200000.0ns 1.089115858078003V 181240000.0ns 1.089115858078003V 181720000.0ns 1.089115858078003V 181760000.0ns 1.089115858078003V 182480000.0ns 1.089115858078003V 182520000.0ns 1.089115858078003V 183000000.0ns 1.089115858078003V 183040000.0ns 1.089115858078003V 183760000.0ns 1.089115858078003V 183800000.0ns 0V 184280000.0ns 0V 184320000.0ns 0.17285370826721191V 185040000.0ns 0.17285370826721191V 185080000.0ns 0.17285370826721191V 185560000.0ns 0.17285370826721191V 185600000.0ns 0.17285370826721191V 186320000.0ns 0.17285370826721191V 186360000.0ns 0.17285370826721191V 186840000.0ns 0.17285370826721191V 186880000.0ns 0.17285370826721191V 187600000.0ns 0.17285370826721191V 187640000.0ns 0V 188120000.0ns 0V 188160000.0ns 0.9819788932800293V 188880000.0ns 0.9819788932800293V 188920000.0ns 0.9819788932800293V 189400000.0ns 0.9819788932800293V 189440000.0ns 0.9819788932800293V 190160000.0ns 0.9819788932800293V 190200000.0ns 0.9819788932800293V 190680000.0ns 0.9819788932800293V 190720000.0ns 0.9819788932800293V 191440000.0ns 0.9819788932800293V 191480000.0ns 0V 191960000.0ns 0V 192000000.0ns 1.9494420289993286V 192720000.0ns 1.9494420289993286V 192760000.0ns 1.9494420289993286V 193240000.0ns 1.9494420289993286V 193280000.0ns 1.9494420289993286V 194000000.0ns 1.9494420289993286V 194040000.0ns 1.9494420289993286V 194520000.0ns 1.9494420289993286V 194560000.0ns 1.9494420289993286V 195280000.0ns 1.9494420289993286V 195320000.0ns 0V 195800000.0ns 0V 195840000.0ns 1.3962270021438599V 196560000.0ns 1.3962270021438599V 196600000.0ns 1.3962270021438599V 197080000.0ns 1.3962270021438599V 197120000.0ns 1.3962270021438599V 197840000.0ns 1.3962270021438599V 197880000.0ns 1.3962270021438599V 198360000.0ns 1.3962270021438599V 198400000.0ns 1.3962270021438599V 199120000.0ns 1.3962270021438599V 199160000.0ns 0V 199640000.0ns 0V 199680000.0ns 1.7114460468292236V 200400000.0ns 1.7114460468292236V 200440000.0ns 1.7114460468292236V 200920000.0ns 1.7114460468292236V 200960000.0ns 1.7114460468292236V 201680000.0ns 1.7114460468292236V 201720000.0ns 1.7114460468292236V 202200000.0ns 1.7114460468292236V 202240000.0ns 1.7114460468292236V 202960000.0ns 1.7114460468292236V 203000000.0ns 0V 203480000.0ns 0V 203520000.0ns 0.9994106292724609V 204240000.0ns 0.9994106292724609V 204280000.0ns 0.9994106292724609V 204760000.0ns 0.9994106292724609V 204800000.0ns 0.9994106292724609V 205520000.0ns 0.9994106292724609V 205560000.0ns 0.9994106292724609V 206040000.0ns 0.9994106292724609V 206080000.0ns 0.9994106292724609V 206800000.0ns 0.9994106292724609V 206840000.0ns 0V 207320000.0ns 0V 207360000.0ns 0.8416277170181274V 208080000.0ns 0.8416277170181274V 208120000.0ns 0.8416277170181274V 208600000.0ns 0.8416277170181274V 208640000.0ns 0.8416277170181274V 209360000.0ns 0.8416277170181274V 209400000.0ns 0.8416277170181274V 209880000.0ns 0.8416277170181274V 209920000.0ns 0.8416277170181274V 210640000.0ns 0.8416277170181274V 210680000.0ns 0V 211160000.0ns 0V 211200000.0ns 1.733735203742981V 211920000.0ns 1.733735203742981V 211960000.0ns 1.733735203742981V 212440000.0ns 1.733735203742981V 212480000.0ns 1.733735203742981V 213200000.0ns 1.733735203742981V 213240000.0ns 1.733735203742981V 213720000.0ns 1.733735203742981V 213760000.0ns 1.733735203742981V 214480000.0ns 1.733735203742981V 214520000.0ns 0V 215000000.0ns 0V 215040000.0ns 0.800771951675415V 215760000.0ns 0.800771951675415V 215800000.0ns 0.800771951675415V 216280000.0ns 0.800771951675415V 216320000.0ns 0.800771951675415V 217040000.0ns 0.800771951675415V 217080000.0ns 0.800771951675415V 217560000.0ns 0.800771951675415V 217600000.0ns 0.800771951675415V 218320000.0ns 0.800771951675415V 218360000.0ns 0V 218840000.0ns 0V 218880000.0ns 1.5126961469650269V 219600000.0ns 1.5126961469650269V 219640000.0ns 1.5126961469650269V 220120000.0ns 1.5126961469650269V 220160000.0ns 1.5126961469650269V 220880000.0ns 1.5126961469650269V 220920000.0ns 1.5126961469650269V 221400000.0ns 1.5126961469650269V 221440000.0ns 1.5126961469650269V 222160000.0ns 1.5126961469650269V 222200000.0ns 0V 222680000.0ns 0V 222720000.0ns 1.5969152450561523V 223440000.0ns 1.5969152450561523V 223480000.0ns 1.5969152450561523V 223960000.0ns 1.5969152450561523V 224000000.0ns 1.5969152450561523V 224720000.0ns 1.5969152450561523V 224760000.0ns 1.5969152450561523V 225240000.0ns 1.5969152450561523V 225280000.0ns 1.5969152450561523V 226000000.0ns 1.5969152450561523V 226040000.0ns 0V 226520000.0ns 0V 226560000.0ns 1.368742823600769V 227280000.0ns 1.368742823600769V 227320000.0ns 1.368742823600769V 227800000.0ns 1.368742823600769V 227840000.0ns 1.368742823600769V 228560000.0ns 1.368742823600769V 228600000.0ns 1.368742823600769V 229080000.0ns 1.368742823600769V 229120000.0ns 1.368742823600769V 229840000.0ns 1.368742823600769V 229880000.0ns 0V 230360000.0ns 0V 230400000.0ns 1.9722808599472046V 231120000.0ns 1.9722808599472046V 231160000.0ns 1.9722808599472046V 231640000.0ns 1.9722808599472046V 231680000.0ns 1.9722808599472046V 232400000.0ns 1.9722808599472046V 232440000.0ns 1.9722808599472046V 232920000.0ns 1.9722808599472046V 232960000.0ns 1.9722808599472046V 233680000.0ns 1.9722808599472046V 233720000.0ns 0V 234200000.0ns 0V 234240000.0ns 0.5916706323623657V 234960000.0ns 0.5916706323623657V 235000000.0ns 0.5916706323623657V 235480000.0ns 0.5916706323623657V 235520000.0ns 0.5916706323623657V 236240000.0ns 0.5916706323623657V 236280000.0ns 0.5916706323623657V 236760000.0ns 0.5916706323623657V 236800000.0ns 0.5916706323623657V 237520000.0ns 0.5916706323623657V 237560000.0ns 0V 238040000.0ns 0V 238080000.0ns 0.7326819896697998V 238800000.0ns 0.7326819896697998V 238840000.0ns 0.7326819896697998V 239320000.0ns 0.7326819896697998V 239360000.0ns 0.7326819896697998V 240080000.0ns 0.7326819896697998V 240120000.0ns 0.7326819896697998V 240600000.0ns 0.7326819896697998V 240640000.0ns 0.7326819896697998V 241360000.0ns 0.7326819896697998V 241400000.0ns 0V 241880000.0ns 0V 241920000.0ns 0.1870344877243042V 242640000.0ns 0.1870344877243042V 242680000.0ns 0.1870344877243042V 243160000.0ns 0.1870344877243042V 243200000.0ns 0.1870344877243042V 243920000.0ns 0.1870344877243042V 243960000.0ns 0.1870344877243042V 244440000.0ns 0.1870344877243042V 244480000.0ns 0.1870344877243042V 245200000.0ns 0.1870344877243042V 245240000.0ns 0V 245720000.0ns 0V 245760000.0ns 0.4935530424118042V 246480000.0ns 0.4935530424118042V 246520000.0ns 0.4935530424118042V 247000000.0ns 0.4935530424118042V 247040000.0ns 0.4935530424118042V 247760000.0ns 0.4935530424118042V 247800000.0ns 0.4935530424118042V 248280000.0ns 0.4935530424118042V 248320000.0ns 0.4935530424118042V 249040000.0ns 0.4935530424118042V 249080000.0ns 0V 249560000.0ns 0V 249600000.0ns 0.11461138725280762V 250320000.0ns 0.11461138725280762V 250360000.0ns 0.11461138725280762V 250840000.0ns 0.11461138725280762V 250880000.0ns 0.11461138725280762V 251600000.0ns 0.11461138725280762V 251640000.0ns 0.11461138725280762V 252120000.0ns 0.11461138725280762V 252160000.0ns 0.11461138725280762V 252880000.0ns 0.11461138725280762V 252920000.0ns 0V 253400000.0ns 0V 253440000.0ns 0.7956382036209106V 254160000.0ns 0.7956382036209106V 254200000.0ns 0.7956382036209106V 254680000.0ns 0.7956382036209106V 254720000.0ns 0.7956382036209106V 255440000.0ns 0.7956382036209106V 255480000.0ns 0.7956382036209106V 255960000.0ns 0.7956382036209106V 256000000.0ns 0.7956382036209106V 256720000.0ns 0.7956382036209106V 256760000.0ns 0V 257240000.0ns 0V 257280000.0ns 1.3353161811828613V 258000000.0ns 1.3353161811828613V 258040000.0ns 1.3353161811828613V 258520000.0ns 1.3353161811828613V 258560000.0ns 1.3353161811828613V 259280000.0ns 1.3353161811828613V 259320000.0ns 1.3353161811828613V 259800000.0ns 1.3353161811828613V 259840000.0ns 1.3353161811828613V 260560000.0ns 1.3353161811828613V 260600000.0ns 0V 261080000.0ns 0V 261120000.0ns 0.07631838321685791V 261840000.0ns 0.07631838321685791V 261880000.0ns 0.07631838321685791V 262360000.0ns 0.07631838321685791V 262400000.0ns 0.07631838321685791V 263120000.0ns 0.07631838321685791V 263160000.0ns 0.07631838321685791V 263640000.0ns 0.07631838321685791V 263680000.0ns 0.07631838321685791V 264400000.0ns 0.07631838321685791V 264440000.0ns 0V 264920000.0ns 0V 264960000.0ns 1.16324782371521V 265680000.0ns 1.16324782371521V 265720000.0ns 1.16324782371521V 266200000.0ns 1.16324782371521V 266240000.0ns 1.16324782371521V 266960000.0ns 1.16324782371521V 267000000.0ns 1.16324782371521V 267480000.0ns 1.16324782371521V 267520000.0ns 1.16324782371521V 268240000.0ns 1.16324782371521V 268280000.0ns 0V 268760000.0ns 0V 268800000.0ns 1.3486560583114624V 269520000.0ns 1.3486560583114624V 269560000.0ns 1.3486560583114624V 270040000.0ns 1.3486560583114624V 270080000.0ns 1.3486560583114624V 270800000.0ns 1.3486560583114624V 270840000.0ns 1.3486560583114624V 271320000.0ns 1.3486560583114624V 271360000.0ns 1.3486560583114624V 272080000.0ns 1.3486560583114624V 272120000.0ns 0V 272600000.0ns 0V 272640000.0ns 0.45393896102905273V 273360000.0ns 0.45393896102905273V 273400000.0ns 0.45393896102905273V 273880000.0ns 0.45393896102905273V 273920000.0ns 0.45393896102905273V 274640000.0ns 0.45393896102905273V 274680000.0ns 0.45393896102905273V 275160000.0ns 0.45393896102905273V 275200000.0ns 0.45393896102905273V 275920000.0ns 0.45393896102905273V 275960000.0ns 0V 276440000.0ns 0V 276480000.0ns 0.7213983535766602V 277200000.0ns 0.7213983535766602V 277240000.0ns 0.7213983535766602V 277720000.0ns 0.7213983535766602V 277760000.0ns 0.7213983535766602V 278480000.0ns 0.7213983535766602V 278520000.0ns 0.7213983535766602V 279000000.0ns 0.7213983535766602V 279040000.0ns 0.7213983535766602V 279760000.0ns 0.7213983535766602V 279800000.0ns 0V 280280000.0ns 0V 280320000.0ns 1.8880258798599243V 281040000.0ns 1.8880258798599243V 281080000.0ns 1.8880258798599243V 281560000.0ns 1.8880258798599243V 281600000.0ns 1.8880258798599243V 282320000.0ns 1.8880258798599243V 282360000.0ns 1.8880258798599243V 282840000.0ns 1.8880258798599243V 282880000.0ns 1.8880258798599243V 283600000.0ns 1.8880258798599243V 283640000.0ns 0V 284120000.0ns 0V 284160000.0ns 0.4708671569824219V 284880000.0ns 0.4708671569824219V 284920000.0ns 0.4708671569824219V 285400000.0ns 0.4708671569824219V 285440000.0ns 0.4708671569824219V 286160000.0ns 0.4708671569824219V 286200000.0ns 0.4708671569824219V 286680000.0ns 0.4708671569824219V 286720000.0ns 0.4708671569824219V 287440000.0ns 0.4708671569824219V 287480000.0ns 0V 287960000.0ns 0V 288000000.0ns 0.9713476896286011V 288720000.0ns 0.9713476896286011V 288760000.0ns 0.9713476896286011V 289240000.0ns 0.9713476896286011V 289280000.0ns 0.9713476896286011V 290000000.0ns 0.9713476896286011V 290040000.0ns 0.9713476896286011V 290520000.0ns 0.9713476896286011V 290560000.0ns 0.9713476896286011V 291280000.0ns 0.9713476896286011V 291320000.0ns 0V 291800000.0ns 0V 291840000.0ns 1.0944520235061646V 292560000.0ns 1.0944520235061646V 292600000.0ns 1.0944520235061646V 293080000.0ns 1.0944520235061646V 293120000.0ns 1.0944520235061646V 293840000.0ns 1.0944520235061646V 293880000.0ns 1.0944520235061646V 294360000.0ns 1.0944520235061646V 294400000.0ns 1.0944520235061646V 295120000.0ns 1.0944520235061646V 295160000.0ns 0V 295640000.0ns 0V 295680000.0ns 1.2067028284072876V 296400000.0ns 1.2067028284072876V 296440000.0ns 1.2067028284072876V 296920000.0ns 1.2067028284072876V 296960000.0ns 1.2067028284072876V 297680000.0ns 1.2067028284072876V 297720000.0ns 1.2067028284072876V 298200000.0ns 1.2067028284072876V 298240000.0ns 1.2067028284072876V 298960000.0ns 1.2067028284072876V 299000000.0ns 0V 299480000.0ns 0V 299520000.0ns 1.9784232378005981V 300240000.0ns 1.9784232378005981V 300280000.0ns 1.9784232378005981V 300760000.0ns 1.9784232378005981V 300800000.0ns 1.9784232378005981V 301520000.0ns 1.9784232378005981V 301560000.0ns 1.9784232378005981V 302040000.0ns 1.9784232378005981V 302080000.0ns 1.9784232378005981V 302800000.0ns 1.9784232378005981V 302840000.0ns 0V 303320000.0ns 0V 303360000.0ns 0.8933771848678589V 304080000.0ns 0.8933771848678589V 304120000.0ns 0.8933771848678589V 304600000.0ns 0.8933771848678589V 304640000.0ns 0.8933771848678589V 305360000.0ns 0.8933771848678589V 305400000.0ns 0.8933771848678589V 305880000.0ns 0.8933771848678589V 305920000.0ns 0.8933771848678589V 306640000.0ns 0.8933771848678589V 306680000.0ns 0V 307160000.0ns 0V 307200000.0ns 1.5887188911437988V 307920000.0ns 1.5887188911437988V 307960000.0ns 1.5887188911437988V 308440000.0ns 1.5887188911437988V 308480000.0ns 1.5887188911437988V 309200000.0ns 1.5887188911437988V 309240000.0ns 1.5887188911437988V 309720000.0ns 1.5887188911437988V 309760000.0ns 1.5887188911437988V 310480000.0ns 1.5887188911437988V 310520000.0ns 0V 311000000.0ns 0V 311040000.0ns 1.588065505027771V 311760000.0ns 1.588065505027771V 311800000.0ns 1.588065505027771V 312280000.0ns 1.588065505027771V 312320000.0ns 1.588065505027771V 313040000.0ns 1.588065505027771V 313080000.0ns 1.588065505027771V 313560000.0ns 1.588065505027771V 313600000.0ns 1.588065505027771V 314320000.0ns 1.588065505027771V 314360000.0ns 0V 314840000.0ns 0V 314880000.0ns 1.192320466041565V 315600000.0ns 1.192320466041565V 315640000.0ns 1.192320466041565V 316120000.0ns 1.192320466041565V 316160000.0ns 1.192320466041565V 316880000.0ns 1.192320466041565V 316920000.0ns 1.192320466041565V 317400000.0ns 1.192320466041565V 317440000.0ns 1.192320466041565V 318160000.0ns 1.192320466041565V 318200000.0ns 0V 318680000.0ns 0V 318720000.0ns 0.7604736089706421V 319440000.0ns 0.7604736089706421V 319480000.0ns 0.7604736089706421V 319960000.0ns 0.7604736089706421V 320000000.0ns 0.7604736089706421V 320720000.0ns 0.7604736089706421V 320760000.0ns 0.7604736089706421V 321240000.0ns 0.7604736089706421V 321280000.0ns 0.7604736089706421V 322000000.0ns 0.7604736089706421V 322040000.0ns 0V 322520000.0ns 0V 322560000.0ns 1.1501935720443726V 323280000.0ns 1.1501935720443726V 323320000.0ns 1.1501935720443726V 323800000.0ns 1.1501935720443726V 323840000.0ns 1.1501935720443726V 324560000.0ns 1.1501935720443726V 324600000.0ns 1.1501935720443726V 325080000.0ns 1.1501935720443726V 325120000.0ns 1.1501935720443726V 325840000.0ns 1.1501935720443726V 325880000.0ns 0V 326360000.0ns 0V 326400000.0ns 0.7045114040374756V 327120000.0ns 0.7045114040374756V 327160000.0ns 0.7045114040374756V 327640000.0ns 0.7045114040374756V 327680000.0ns 0.7045114040374756V 328400000.0ns 0.7045114040374756V 328440000.0ns 0.7045114040374756V 328920000.0ns 0.7045114040374756V 328960000.0ns 0.7045114040374756V 329680000.0ns 0.7045114040374756V 329720000.0ns 0V 330200000.0ns 0V 330240000.0ns 0.4002110958099365V 330960000.0ns 0.4002110958099365V 331000000.0ns 0.4002110958099365V 331480000.0ns 0.4002110958099365V 331520000.0ns 0.4002110958099365V 332240000.0ns 0.4002110958099365V 332280000.0ns 0.4002110958099365V 332760000.0ns 0.4002110958099365V 332800000.0ns 0.4002110958099365V 333520000.0ns 0.4002110958099365V 333560000.0ns 0V 334040000.0ns 0V 334080000.0ns 1.2367199659347534V 334800000.0ns 1.2367199659347534V 334840000.0ns 1.2367199659347534V 335320000.0ns 1.2367199659347534V 335360000.0ns 1.2367199659347534V 336080000.0ns 1.2367199659347534V 336120000.0ns 1.2367199659347534V 336600000.0ns 1.2367199659347534V 336640000.0ns 1.2367199659347534V 337360000.0ns 1.2367199659347534V 337400000.0ns 0V 337880000.0ns 0V 337920000.0ns 1.941900372505188V 338640000.0ns 1.941900372505188V 338680000.0ns 1.941900372505188V 339160000.0ns 1.941900372505188V 339200000.0ns 1.941900372505188V 339920000.0ns 1.941900372505188V 339960000.0ns 1.941900372505188V 340440000.0ns 1.941900372505188V 340480000.0ns 1.941900372505188V 341200000.0ns 1.941900372505188V 341240000.0ns 0V 341720000.0ns 0V 341760000.0ns 0.5684245824813843V 342480000.0ns 0.5684245824813843V 342520000.0ns 0.5684245824813843V 343000000.0ns 0.5684245824813843V 343040000.0ns 0.5684245824813843V 343760000.0ns 0.5684245824813843V 343800000.0ns 0.5684245824813843V 344280000.0ns 0.5684245824813843V 344320000.0ns 0.5684245824813843V 345040000.0ns 0.5684245824813843V 345080000.0ns 0V 345560000.0ns 0V 345600000.0ns 0.33742809295654297V 346320000.0ns 0.33742809295654297V 346360000.0ns 0.33742809295654297V 346840000.0ns 0.33742809295654297V 346880000.0ns 0.33742809295654297V 347600000.0ns 0.33742809295654297V 347640000.0ns 0.33742809295654297V 348120000.0ns 0.33742809295654297V 348160000.0ns 0.33742809295654297V 348880000.0ns 0.33742809295654297V 348920000.0ns 0V 349400000.0ns 0V 349440000.0ns 1.1796358823776245V 350160000.0ns 1.1796358823776245V 350200000.0ns 1.1796358823776245V 350680000.0ns 1.1796358823776245V 350720000.0ns 1.1796358823776245V 351440000.0ns 1.1796358823776245V 351480000.0ns 1.1796358823776245V 351960000.0ns 1.1796358823776245V 352000000.0ns 1.1796358823776245V 352720000.0ns 1.1796358823776245V 352760000.0ns 0V 353240000.0ns 0V 353280000.0ns 0.36788618564605713V 354000000.0ns 0.36788618564605713V 354040000.0ns 0.36788618564605713V 354520000.0ns 0.36788618564605713V 354560000.0ns 0.36788618564605713V 355280000.0ns 0.36788618564605713V 355320000.0ns 0.36788618564605713V 355800000.0ns 0.36788618564605713V 355840000.0ns 0.36788618564605713V 356560000.0ns 0.36788618564605713V 356600000.0ns 0V 357080000.0ns 0V 357120000.0ns 1.4921669960021973V 357840000.0ns 1.4921669960021973V 357880000.0ns 1.4921669960021973V 358360000.0ns 1.4921669960021973V 358400000.0ns 1.4921669960021973V 359120000.0ns 1.4921669960021973V 359160000.0ns 1.4921669960021973V 359640000.0ns 1.4921669960021973V 359680000.0ns 1.4921669960021973V 360400000.0ns 1.4921669960021973V 360440000.0ns 0V 360920000.0ns 0V 360960000.0ns 1.4613587856292725V 361680000.0ns 1.4613587856292725V 361720000.0ns 1.4613587856292725V 362200000.0ns 1.4613587856292725V 362240000.0ns 1.4613587856292725V 362960000.0ns 1.4613587856292725V 363000000.0ns 1.4613587856292725V 363480000.0ns 1.4613587856292725V 363520000.0ns 1.4613587856292725V 364240000.0ns 1.4613587856292725V 364280000.0ns 0V 364760000.0ns 0V 364800000.0ns 1.0565704107284546V 365520000.0ns 1.0565704107284546V 365560000.0ns 1.0565704107284546V 366040000.0ns 1.0565704107284546V 366080000.0ns 1.0565704107284546V 366800000.0ns 1.0565704107284546V 366840000.0ns 1.0565704107284546V 367320000.0ns 1.0565704107284546V 367360000.0ns 1.0565704107284546V 368080000.0ns 1.0565704107284546V 368120000.0ns 0V 368600000.0ns 0V 368640000.0ns 0.38741743564605713V 369360000.0ns 0.38741743564605713V 369400000.0ns 0.38741743564605713V 369880000.0ns 0.38741743564605713V 369920000.0ns 0.38741743564605713V 370640000.0ns 0.38741743564605713V 370680000.0ns 0.38741743564605713V 371160000.0ns 0.38741743564605713V 371200000.0ns 0.38741743564605713V 371920000.0ns 0.38741743564605713V 371960000.0ns 0V 372440000.0ns 0V 372480000.0ns 0.8422540426254272V 373200000.0ns 0.8422540426254272V 373240000.0ns 0.8422540426254272V 373720000.0ns 0.8422540426254272V 373760000.0ns 0.8422540426254272V 374480000.0ns 0.8422540426254272V 374520000.0ns 0.8422540426254272V 375000000.0ns 0.8422540426254272V 375040000.0ns 0.8422540426254272V 375760000.0ns 0.8422540426254272V 375800000.0ns 0V 376280000.0ns 0V 376320000.0ns 0.034389376640319824V 377040000.0ns 0.034389376640319824V 377080000.0ns 0.034389376640319824V 377560000.0ns 0.034389376640319824V 377600000.0ns 0.034389376640319824V 378320000.0ns 0.034389376640319824V 378360000.0ns 0.034389376640319824V 378840000.0ns 0.034389376640319824V 378880000.0ns 0.034389376640319824V 379600000.0ns 0.034389376640319824V 379640000.0ns 0V 380120000.0ns 0V 380160000.0ns 0.8860955238342285V 380880000.0ns 0.8860955238342285V 380920000.0ns 0.8860955238342285V 381400000.0ns 0.8860955238342285V 381440000.0ns 0.8860955238342285V 382160000.0ns 0.8860955238342285V 382200000.0ns 0.8860955238342285V 382680000.0ns 0.8860955238342285V 382720000.0ns 0.8860955238342285V 383440000.0ns 0.8860955238342285V 383480000.0ns 0V 383960000.0ns 0V 384000000.0ns 0.7267136573791504V 384720000.0ns 0.7267136573791504V 384760000.0ns 0.7267136573791504V 385240000.0ns 0.7267136573791504V 385280000.0ns 0.7267136573791504V 386000000.0ns 0.7267136573791504V 386040000.0ns 0.7267136573791504V 386520000.0ns 0.7267136573791504V 386560000.0ns 0.7267136573791504V 387280000.0ns 0.7267136573791504V 387320000.0ns 0V 387800000.0ns 0V 387840000.0ns 0.3769960403442383V 388560000.0ns 0.3769960403442383V 388600000.0ns 0.3769960403442383V 389080000.0ns 0.3769960403442383V 389120000.0ns 0.3769960403442383V 389840000.0ns 0.3769960403442383V 389880000.0ns 0.3769960403442383V 390360000.0ns 0.3769960403442383V 390400000.0ns 0.3769960403442383V 391120000.0ns 0.3769960403442383V 391160000.0ns 0V)
VX_2 X_2 0 PWL(0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 2.0V 8400000.0ns 2.0V 8440000.0ns 2.0V 8920000.0ns 2.0V 8960000.0ns 2.0V 9680000.0ns 2.0V 9720000.0ns 2.0V 10200000.0ns 2.0V 10240000.0ns 2.0V 10960000.0ns 2.0V 11000000.0ns 0V 11480000.0ns 0V 11520000.0ns 2.0V 12240000.0ns 2.0V 12280000.0ns 2.0V 12760000.0ns 2.0V 12800000.0ns 2.0V 13520000.0ns 2.0V 13560000.0ns 2.0V 14040000.0ns 2.0V 14080000.0ns 2.0V 14800000.0ns 2.0V 14840000.0ns 0V 15320000.0ns 0V 15360000.0ns 2.0V 16080000.0ns 2.0V 16120000.0ns 2.0V 16600000.0ns 2.0V 16640000.0ns 2.0V 17360000.0ns 2.0V 17400000.0ns 2.0V 17880000.0ns 2.0V 17920000.0ns 2.0V 18640000.0ns 2.0V 18680000.0ns 0V 19160000.0ns 0V 19200000.0ns 2.0V 19920000.0ns 2.0V 19960000.0ns 2.0V 20440000.0ns 2.0V 20480000.0ns 2.0V 21200000.0ns 2.0V 21240000.0ns 2.0V 21720000.0ns 2.0V 21760000.0ns 2.0V 22480000.0ns 2.0V 22520000.0ns 0V 23000000.0ns 0V 23040000.0ns 2.0V 23760000.0ns 2.0V 23800000.0ns 2.0V 24280000.0ns 2.0V 24320000.0ns 2.0V 25040000.0ns 2.0V 25080000.0ns 2.0V 25560000.0ns 2.0V 25600000.0ns 2.0V 26320000.0ns 2.0V 26360000.0ns 0V 26840000.0ns 0V 26880000.0ns 2.0V 27600000.0ns 2.0V 27640000.0ns 2.0V 28120000.0ns 2.0V 28160000.0ns 2.0V 28880000.0ns 2.0V 28920000.0ns 2.0V 29400000.0ns 2.0V 29440000.0ns 2.0V 30160000.0ns 2.0V 30200000.0ns 0V 30680000.0ns 0V 30720000.0ns 2.0V 31440000.0ns 2.0V 31480000.0ns 2.0V 31960000.0ns 2.0V 32000000.0ns 2.0V 32720000.0ns 2.0V 32760000.0ns 2.0V 33240000.0ns 2.0V 33280000.0ns 2.0V 34000000.0ns 2.0V 34040000.0ns 0V 34520000.0ns 0V 34560000.0ns 2.0V 35280000.0ns 2.0V 35320000.0ns 2.0V 35800000.0ns 2.0V 35840000.0ns 2.0V 36560000.0ns 2.0V 36600000.0ns 2.0V 37080000.0ns 2.0V 37120000.0ns 2.0V 37840000.0ns 2.0V 37880000.0ns 0V 38360000.0ns 0V 38400000.0ns 2.0V 39120000.0ns 2.0V 39160000.0ns 2.0V 39640000.0ns 2.0V 39680000.0ns 2.0V 40400000.0ns 2.0V 40440000.0ns 2.0V 40920000.0ns 2.0V 40960000.0ns 2.0V 41680000.0ns 2.0V 41720000.0ns 0V 42200000.0ns 0V 42240000.0ns 2.0V 42960000.0ns 2.0V 43000000.0ns 2.0V 43480000.0ns 2.0V 43520000.0ns 2.0V 44240000.0ns 2.0V 44280000.0ns 2.0V 44760000.0ns 2.0V 44800000.0ns 2.0V 45520000.0ns 2.0V 45560000.0ns 0V 46040000.0ns 0V 46080000.0ns 2.0V 46800000.0ns 2.0V 46840000.0ns 2.0V 47320000.0ns 2.0V 47360000.0ns 2.0V 48080000.0ns 2.0V 48120000.0ns 2.0V 48600000.0ns 2.0V 48640000.0ns 2.0V 49360000.0ns 2.0V 49400000.0ns 0V 49880000.0ns 0V 49920000.0ns 2.0V 50640000.0ns 2.0V 50680000.0ns 2.0V 51160000.0ns 2.0V 51200000.0ns 2.0V 51920000.0ns 2.0V 51960000.0ns 2.0V 52440000.0ns 2.0V 52480000.0ns 2.0V 53200000.0ns 2.0V 53240000.0ns 0V 53720000.0ns 0V 53760000.0ns 2.0V 54480000.0ns 2.0V 54520000.0ns 2.0V 55000000.0ns 2.0V 55040000.0ns 2.0V 55760000.0ns 2.0V 55800000.0ns 2.0V 56280000.0ns 2.0V 56320000.0ns 2.0V 57040000.0ns 2.0V 57080000.0ns 0V 57560000.0ns 0V 57600000.0ns 2.0V 58320000.0ns 2.0V 58360000.0ns 2.0V 58840000.0ns 2.0V 58880000.0ns 2.0V 59600000.0ns 2.0V 59640000.0ns 2.0V 60120000.0ns 2.0V 60160000.0ns 2.0V 60880000.0ns 2.0V 60920000.0ns 0V 61400000.0ns 0V 61440000.0ns 2.0V 62160000.0ns 2.0V 62200000.0ns 2.0V 62680000.0ns 2.0V 62720000.0ns 2.0V 63440000.0ns 2.0V 63480000.0ns 2.0V 63960000.0ns 2.0V 64000000.0ns 2.0V 64720000.0ns 2.0V 64760000.0ns 0V 65240000.0ns 0V 65280000.0ns 2.0V 66000000.0ns 2.0V 66040000.0ns 2.0V 66520000.0ns 2.0V 66560000.0ns 2.0V 67280000.0ns 2.0V 67320000.0ns 2.0V 67800000.0ns 2.0V 67840000.0ns 2.0V 68560000.0ns 2.0V 68600000.0ns 0V 69080000.0ns 0V 69120000.0ns 2.0V 69840000.0ns 2.0V 69880000.0ns 2.0V 70360000.0ns 2.0V 70400000.0ns 2.0V 71120000.0ns 2.0V 71160000.0ns 2.0V 71640000.0ns 2.0V 71680000.0ns 2.0V 72400000.0ns 2.0V 72440000.0ns 0V 72920000.0ns 0V 72960000.0ns 2.0V 73680000.0ns 2.0V 73720000.0ns 2.0V 74200000.0ns 2.0V 74240000.0ns 2.0V 74960000.0ns 2.0V 75000000.0ns 2.0V 75480000.0ns 2.0V 75520000.0ns 2.0V 76240000.0ns 2.0V 76280000.0ns 0V 76760000.0ns 0V 76800000.0ns 2.0V 77520000.0ns 2.0V 77560000.0ns 2.0V 78040000.0ns 2.0V 78080000.0ns 2.0V 78800000.0ns 2.0V 78840000.0ns 2.0V 79320000.0ns 2.0V 79360000.0ns 2.0V 80080000.0ns 2.0V 80120000.0ns 0V 80600000.0ns 0V 80640000.0ns 2.0V 81360000.0ns 2.0V 81400000.0ns 2.0V 81880000.0ns 2.0V 81920000.0ns 2.0V 82640000.0ns 2.0V 82680000.0ns 2.0V 83160000.0ns 2.0V 83200000.0ns 2.0V 83920000.0ns 2.0V 83960000.0ns 0V 84440000.0ns 0V 84480000.0ns 2.0V 85200000.0ns 2.0V 85240000.0ns 2.0V 85720000.0ns 2.0V 85760000.0ns 2.0V 86480000.0ns 2.0V 86520000.0ns 2.0V 87000000.0ns 2.0V 87040000.0ns 2.0V 87760000.0ns 2.0V 87800000.0ns 0V 88280000.0ns 0V 88320000.0ns 2.0V 89040000.0ns 2.0V 89080000.0ns 2.0V 89560000.0ns 2.0V 89600000.0ns 2.0V 90320000.0ns 2.0V 90360000.0ns 2.0V 90840000.0ns 2.0V 90880000.0ns 2.0V 91600000.0ns 2.0V 91640000.0ns 0V 92120000.0ns 0V 92160000.0ns 2.0V 92880000.0ns 2.0V 92920000.0ns 2.0V 93400000.0ns 2.0V 93440000.0ns 2.0V 94160000.0ns 2.0V 94200000.0ns 2.0V 94680000.0ns 2.0V 94720000.0ns 2.0V 95440000.0ns 2.0V 95480000.0ns 0V 95960000.0ns 0V 96000000.0ns 2.0V 96720000.0ns 2.0V 96760000.0ns 2.0V 97240000.0ns 2.0V 97280000.0ns 2.0V 98000000.0ns 2.0V 98040000.0ns 2.0V 98520000.0ns 2.0V 98560000.0ns 2.0V 99280000.0ns 2.0V 99320000.0ns 0V 99800000.0ns 0V 99840000.0ns 2.0V 100560000.0ns 2.0V 100600000.0ns 2.0V 101080000.0ns 2.0V 101120000.0ns 2.0V 101840000.0ns 2.0V 101880000.0ns 2.0V 102360000.0ns 2.0V 102400000.0ns 2.0V 103120000.0ns 2.0V 103160000.0ns 0V 103640000.0ns 0V 103680000.0ns 2.0V 104400000.0ns 2.0V 104440000.0ns 2.0V 104920000.0ns 2.0V 104960000.0ns 2.0V 105680000.0ns 2.0V 105720000.0ns 2.0V 106200000.0ns 2.0V 106240000.0ns 2.0V 106960000.0ns 2.0V 107000000.0ns 0V 107480000.0ns 0V 107520000.0ns 2.0V 108240000.0ns 2.0V 108280000.0ns 2.0V 108760000.0ns 2.0V 108800000.0ns 2.0V 109520000.0ns 2.0V 109560000.0ns 2.0V 110040000.0ns 2.0V 110080000.0ns 2.0V 110800000.0ns 2.0V 110840000.0ns 0V 111320000.0ns 0V 111360000.0ns 2.0V 112080000.0ns 2.0V 112120000.0ns 2.0V 112600000.0ns 2.0V 112640000.0ns 2.0V 113360000.0ns 2.0V 113400000.0ns 2.0V 113880000.0ns 2.0V 113920000.0ns 2.0V 114640000.0ns 2.0V 114680000.0ns 0V 115160000.0ns 0V 115200000.0ns 2.0V 115920000.0ns 2.0V 115960000.0ns 2.0V 116440000.0ns 2.0V 116480000.0ns 2.0V 117200000.0ns 2.0V 117240000.0ns 2.0V 117720000.0ns 2.0V 117760000.0ns 2.0V 118480000.0ns 2.0V 118520000.0ns 0V 119000000.0ns 0V 119040000.0ns 2.0V 119760000.0ns 2.0V 119800000.0ns 2.0V 120280000.0ns 2.0V 120320000.0ns 2.0V 121040000.0ns 2.0V 121080000.0ns 2.0V 121560000.0ns 2.0V 121600000.0ns 2.0V 122320000.0ns 2.0V 122360000.0ns 0V 122840000.0ns 0V 122880000.0ns 2.0V 123600000.0ns 2.0V 123640000.0ns 2.0V 124120000.0ns 2.0V 124160000.0ns 2.0V 124880000.0ns 2.0V 124920000.0ns 2.0V 125400000.0ns 2.0V 125440000.0ns 2.0V 126160000.0ns 2.0V 126200000.0ns 0V 126680000.0ns 0V 126720000.0ns 2.0V 127440000.0ns 2.0V 127480000.0ns 2.0V 127960000.0ns 2.0V 128000000.0ns 2.0V 128720000.0ns 2.0V 128760000.0ns 2.0V 129240000.0ns 2.0V 129280000.0ns 2.0V 130000000.0ns 2.0V 130040000.0ns 0V 130520000.0ns 0V 130560000.0ns 2.0V 131280000.0ns 2.0V 131320000.0ns 2.0V 131800000.0ns 2.0V 131840000.0ns 2.0V 132560000.0ns 2.0V 132600000.0ns 2.0V 133080000.0ns 2.0V 133120000.0ns 2.0V 133840000.0ns 2.0V 133880000.0ns 0V 134360000.0ns 0V 134400000.0ns 2.0V 135120000.0ns 2.0V 135160000.0ns 2.0V 135640000.0ns 2.0V 135680000.0ns 2.0V 136400000.0ns 2.0V 136440000.0ns 2.0V 136920000.0ns 2.0V 136960000.0ns 2.0V 137680000.0ns 2.0V 137720000.0ns 0V 138200000.0ns 0V 138240000.0ns 2.0V 138960000.0ns 2.0V 139000000.0ns 2.0V 139480000.0ns 2.0V 139520000.0ns 2.0V 140240000.0ns 2.0V 140280000.0ns 2.0V 140760000.0ns 2.0V 140800000.0ns 2.0V 141520000.0ns 2.0V 141560000.0ns 0V 142040000.0ns 0V 142080000.0ns 2.0V 142800000.0ns 2.0V 142840000.0ns 2.0V 143320000.0ns 2.0V 143360000.0ns 2.0V 144080000.0ns 2.0V 144120000.0ns 2.0V 144600000.0ns 2.0V 144640000.0ns 2.0V 145360000.0ns 2.0V 145400000.0ns 0V 145880000.0ns 0V 145920000.0ns 2.0V 146640000.0ns 2.0V 146680000.0ns 2.0V 147160000.0ns 2.0V 147200000.0ns 2.0V 147920000.0ns 2.0V 147960000.0ns 2.0V 148440000.0ns 2.0V 148480000.0ns 2.0V 149200000.0ns 2.0V 149240000.0ns 0V 149720000.0ns 0V 149760000.0ns 2.0V 150480000.0ns 2.0V 150520000.0ns 2.0V 151000000.0ns 2.0V 151040000.0ns 2.0V 151760000.0ns 2.0V 151800000.0ns 2.0V 152280000.0ns 2.0V 152320000.0ns 2.0V 153040000.0ns 2.0V 153080000.0ns 0V 153560000.0ns 0V 153600000.0ns 2.0V 154320000.0ns 2.0V 154360000.0ns 2.0V 154840000.0ns 2.0V 154880000.0ns 2.0V 155600000.0ns 2.0V 155640000.0ns 2.0V 156120000.0ns 2.0V 156160000.0ns 2.0V 156880000.0ns 2.0V 156920000.0ns 0V 157400000.0ns 0V 157440000.0ns 2.0V 158160000.0ns 2.0V 158200000.0ns 2.0V 158680000.0ns 2.0V 158720000.0ns 2.0V 159440000.0ns 2.0V 159480000.0ns 2.0V 159960000.0ns 2.0V 160000000.0ns 2.0V 160720000.0ns 2.0V 160760000.0ns 0V 161240000.0ns 0V 161280000.0ns 2.0V 162000000.0ns 2.0V 162040000.0ns 2.0V 162520000.0ns 2.0V 162560000.0ns 2.0V 163280000.0ns 2.0V 163320000.0ns 2.0V 163800000.0ns 2.0V 163840000.0ns 2.0V 164560000.0ns 2.0V 164600000.0ns 0V 165080000.0ns 0V 165120000.0ns 2.0V 165840000.0ns 2.0V 165880000.0ns 2.0V 166360000.0ns 2.0V 166400000.0ns 2.0V 167120000.0ns 2.0V 167160000.0ns 2.0V 167640000.0ns 2.0V 167680000.0ns 2.0V 168400000.0ns 2.0V 168440000.0ns 0V 168920000.0ns 0V 168960000.0ns 2.0V 169680000.0ns 2.0V 169720000.0ns 2.0V 170200000.0ns 2.0V 170240000.0ns 2.0V 170960000.0ns 2.0V 171000000.0ns 2.0V 171480000.0ns 2.0V 171520000.0ns 2.0V 172240000.0ns 2.0V 172280000.0ns 0V 172760000.0ns 0V 172800000.0ns 2.0V 173520000.0ns 2.0V 173560000.0ns 2.0V 174040000.0ns 2.0V 174080000.0ns 2.0V 174800000.0ns 2.0V 174840000.0ns 2.0V 175320000.0ns 2.0V 175360000.0ns 2.0V 176080000.0ns 2.0V 176120000.0ns 0V 176600000.0ns 0V 176640000.0ns 2.0V 177360000.0ns 2.0V 177400000.0ns 2.0V 177880000.0ns 2.0V 177920000.0ns 2.0V 178640000.0ns 2.0V 178680000.0ns 2.0V 179160000.0ns 2.0V 179200000.0ns 2.0V 179920000.0ns 2.0V 179960000.0ns 0V 180440000.0ns 0V 180480000.0ns 2.0V 181200000.0ns 2.0V 181240000.0ns 2.0V 181720000.0ns 2.0V 181760000.0ns 2.0V 182480000.0ns 2.0V 182520000.0ns 2.0V 183000000.0ns 2.0V 183040000.0ns 2.0V 183760000.0ns 2.0V 183800000.0ns 0V 184280000.0ns 0V 184320000.0ns 2.0V 185040000.0ns 2.0V 185080000.0ns 2.0V 185560000.0ns 2.0V 185600000.0ns 2.0V 186320000.0ns 2.0V 186360000.0ns 2.0V 186840000.0ns 2.0V 186880000.0ns 2.0V 187600000.0ns 2.0V 187640000.0ns 0V 188120000.0ns 0V 188160000.0ns 2.0V 188880000.0ns 2.0V 188920000.0ns 2.0V 189400000.0ns 2.0V 189440000.0ns 2.0V 190160000.0ns 2.0V 190200000.0ns 2.0V 190680000.0ns 2.0V 190720000.0ns 2.0V 191440000.0ns 2.0V 191480000.0ns 0V 191960000.0ns 0V 192000000.0ns 2.0V 192720000.0ns 2.0V 192760000.0ns 2.0V 193240000.0ns 2.0V 193280000.0ns 2.0V 194000000.0ns 2.0V 194040000.0ns 2.0V 194520000.0ns 2.0V 194560000.0ns 2.0V 195280000.0ns 2.0V 195320000.0ns 0V 195800000.0ns 0V 195840000.0ns 2.0V 196560000.0ns 2.0V 196600000.0ns 2.0V 197080000.0ns 2.0V 197120000.0ns 2.0V 197840000.0ns 2.0V 197880000.0ns 2.0V 198360000.0ns 2.0V 198400000.0ns 2.0V 199120000.0ns 2.0V 199160000.0ns 0V 199640000.0ns 0V 199680000.0ns 2.0V 200400000.0ns 2.0V 200440000.0ns 2.0V 200920000.0ns 2.0V 200960000.0ns 2.0V 201680000.0ns 2.0V 201720000.0ns 2.0V 202200000.0ns 2.0V 202240000.0ns 2.0V 202960000.0ns 2.0V 203000000.0ns 0V 203480000.0ns 0V 203520000.0ns 2.0V 204240000.0ns 2.0V 204280000.0ns 2.0V 204760000.0ns 2.0V 204800000.0ns 2.0V 205520000.0ns 2.0V 205560000.0ns 2.0V 206040000.0ns 2.0V 206080000.0ns 2.0V 206800000.0ns 2.0V 206840000.0ns 0V 207320000.0ns 0V 207360000.0ns 2.0V 208080000.0ns 2.0V 208120000.0ns 2.0V 208600000.0ns 2.0V 208640000.0ns 2.0V 209360000.0ns 2.0V 209400000.0ns 2.0V 209880000.0ns 2.0V 209920000.0ns 2.0V 210640000.0ns 2.0V 210680000.0ns 0V 211160000.0ns 0V 211200000.0ns 2.0V 211920000.0ns 2.0V 211960000.0ns 2.0V 212440000.0ns 2.0V 212480000.0ns 2.0V 213200000.0ns 2.0V 213240000.0ns 2.0V 213720000.0ns 2.0V 213760000.0ns 2.0V 214480000.0ns 2.0V 214520000.0ns 0V 215000000.0ns 0V 215040000.0ns 2.0V 215760000.0ns 2.0V 215800000.0ns 2.0V 216280000.0ns 2.0V 216320000.0ns 2.0V 217040000.0ns 2.0V 217080000.0ns 2.0V 217560000.0ns 2.0V 217600000.0ns 2.0V 218320000.0ns 2.0V 218360000.0ns 0V 218840000.0ns 0V 218880000.0ns 2.0V 219600000.0ns 2.0V 219640000.0ns 2.0V 220120000.0ns 2.0V 220160000.0ns 2.0V 220880000.0ns 2.0V 220920000.0ns 2.0V 221400000.0ns 2.0V 221440000.0ns 2.0V 222160000.0ns 2.0V 222200000.0ns 0V 222680000.0ns 0V 222720000.0ns 2.0V 223440000.0ns 2.0V 223480000.0ns 2.0V 223960000.0ns 2.0V 224000000.0ns 2.0V 224720000.0ns 2.0V 224760000.0ns 2.0V 225240000.0ns 2.0V 225280000.0ns 2.0V 226000000.0ns 2.0V 226040000.0ns 0V 226520000.0ns 0V 226560000.0ns 2.0V 227280000.0ns 2.0V 227320000.0ns 2.0V 227800000.0ns 2.0V 227840000.0ns 2.0V 228560000.0ns 2.0V 228600000.0ns 2.0V 229080000.0ns 2.0V 229120000.0ns 2.0V 229840000.0ns 2.0V 229880000.0ns 0V 230360000.0ns 0V 230400000.0ns 2.0V 231120000.0ns 2.0V 231160000.0ns 2.0V 231640000.0ns 2.0V 231680000.0ns 2.0V 232400000.0ns 2.0V 232440000.0ns 2.0V 232920000.0ns 2.0V 232960000.0ns 2.0V 233680000.0ns 2.0V 233720000.0ns 0V 234200000.0ns 0V 234240000.0ns 2.0V 234960000.0ns 2.0V 235000000.0ns 2.0V 235480000.0ns 2.0V 235520000.0ns 2.0V 236240000.0ns 2.0V 236280000.0ns 2.0V 236760000.0ns 2.0V 236800000.0ns 2.0V 237520000.0ns 2.0V 237560000.0ns 0V 238040000.0ns 0V 238080000.0ns 2.0V 238800000.0ns 2.0V 238840000.0ns 2.0V 239320000.0ns 2.0V 239360000.0ns 2.0V 240080000.0ns 2.0V 240120000.0ns 2.0V 240600000.0ns 2.0V 240640000.0ns 2.0V 241360000.0ns 2.0V 241400000.0ns 0V 241880000.0ns 0V 241920000.0ns 2.0V 242640000.0ns 2.0V 242680000.0ns 2.0V 243160000.0ns 2.0V 243200000.0ns 2.0V 243920000.0ns 2.0V 243960000.0ns 2.0V 244440000.0ns 2.0V 244480000.0ns 2.0V 245200000.0ns 2.0V 245240000.0ns 0V 245720000.0ns 0V 245760000.0ns 2.0V 246480000.0ns 2.0V 246520000.0ns 2.0V 247000000.0ns 2.0V 247040000.0ns 2.0V 247760000.0ns 2.0V 247800000.0ns 2.0V 248280000.0ns 2.0V 248320000.0ns 2.0V 249040000.0ns 2.0V 249080000.0ns 0V 249560000.0ns 0V 249600000.0ns 2.0V 250320000.0ns 2.0V 250360000.0ns 2.0V 250840000.0ns 2.0V 250880000.0ns 2.0V 251600000.0ns 2.0V 251640000.0ns 2.0V 252120000.0ns 2.0V 252160000.0ns 2.0V 252880000.0ns 2.0V 252920000.0ns 0V 253400000.0ns 0V 253440000.0ns 2.0V 254160000.0ns 2.0V 254200000.0ns 2.0V 254680000.0ns 2.0V 254720000.0ns 2.0V 255440000.0ns 2.0V 255480000.0ns 2.0V 255960000.0ns 2.0V 256000000.0ns 2.0V 256720000.0ns 2.0V 256760000.0ns 0V 257240000.0ns 0V 257280000.0ns 2.0V 258000000.0ns 2.0V 258040000.0ns 2.0V 258520000.0ns 2.0V 258560000.0ns 2.0V 259280000.0ns 2.0V 259320000.0ns 2.0V 259800000.0ns 2.0V 259840000.0ns 2.0V 260560000.0ns 2.0V 260600000.0ns 0V 261080000.0ns 0V 261120000.0ns 2.0V 261840000.0ns 2.0V 261880000.0ns 2.0V 262360000.0ns 2.0V 262400000.0ns 2.0V 263120000.0ns 2.0V 263160000.0ns 2.0V 263640000.0ns 2.0V 263680000.0ns 2.0V 264400000.0ns 2.0V 264440000.0ns 0V 264920000.0ns 0V 264960000.0ns 2.0V 265680000.0ns 2.0V 265720000.0ns 2.0V 266200000.0ns 2.0V 266240000.0ns 2.0V 266960000.0ns 2.0V 267000000.0ns 2.0V 267480000.0ns 2.0V 267520000.0ns 2.0V 268240000.0ns 2.0V 268280000.0ns 0V 268760000.0ns 0V 268800000.0ns 2.0V 269520000.0ns 2.0V 269560000.0ns 2.0V 270040000.0ns 2.0V 270080000.0ns 2.0V 270800000.0ns 2.0V 270840000.0ns 2.0V 271320000.0ns 2.0V 271360000.0ns 2.0V 272080000.0ns 2.0V 272120000.0ns 0V 272600000.0ns 0V 272640000.0ns 2.0V 273360000.0ns 2.0V 273400000.0ns 2.0V 273880000.0ns 2.0V 273920000.0ns 2.0V 274640000.0ns 2.0V 274680000.0ns 2.0V 275160000.0ns 2.0V 275200000.0ns 2.0V 275920000.0ns 2.0V 275960000.0ns 0V 276440000.0ns 0V 276480000.0ns 2.0V 277200000.0ns 2.0V 277240000.0ns 2.0V 277720000.0ns 2.0V 277760000.0ns 2.0V 278480000.0ns 2.0V 278520000.0ns 2.0V 279000000.0ns 2.0V 279040000.0ns 2.0V 279760000.0ns 2.0V 279800000.0ns 0V 280280000.0ns 0V 280320000.0ns 2.0V 281040000.0ns 2.0V 281080000.0ns 2.0V 281560000.0ns 2.0V 281600000.0ns 2.0V 282320000.0ns 2.0V 282360000.0ns 2.0V 282840000.0ns 2.0V 282880000.0ns 2.0V 283600000.0ns 2.0V 283640000.0ns 0V 284120000.0ns 0V 284160000.0ns 2.0V 284880000.0ns 2.0V 284920000.0ns 2.0V 285400000.0ns 2.0V 285440000.0ns 2.0V 286160000.0ns 2.0V 286200000.0ns 2.0V 286680000.0ns 2.0V 286720000.0ns 2.0V 287440000.0ns 2.0V 287480000.0ns 0V 287960000.0ns 0V 288000000.0ns 2.0V 288720000.0ns 2.0V 288760000.0ns 2.0V 289240000.0ns 2.0V 289280000.0ns 2.0V 290000000.0ns 2.0V 290040000.0ns 2.0V 290520000.0ns 2.0V 290560000.0ns 2.0V 291280000.0ns 2.0V 291320000.0ns 0V 291800000.0ns 0V 291840000.0ns 2.0V 292560000.0ns 2.0V 292600000.0ns 2.0V 293080000.0ns 2.0V 293120000.0ns 2.0V 293840000.0ns 2.0V 293880000.0ns 2.0V 294360000.0ns 2.0V 294400000.0ns 2.0V 295120000.0ns 2.0V 295160000.0ns 0V 295640000.0ns 0V 295680000.0ns 2.0V 296400000.0ns 2.0V 296440000.0ns 2.0V 296920000.0ns 2.0V 296960000.0ns 2.0V 297680000.0ns 2.0V 297720000.0ns 2.0V 298200000.0ns 2.0V 298240000.0ns 2.0V 298960000.0ns 2.0V 299000000.0ns 0V 299480000.0ns 0V 299520000.0ns 2.0V 300240000.0ns 2.0V 300280000.0ns 2.0V 300760000.0ns 2.0V 300800000.0ns 2.0V 301520000.0ns 2.0V 301560000.0ns 2.0V 302040000.0ns 2.0V 302080000.0ns 2.0V 302800000.0ns 2.0V 302840000.0ns 0V 303320000.0ns 0V 303360000.0ns 2.0V 304080000.0ns 2.0V 304120000.0ns 2.0V 304600000.0ns 2.0V 304640000.0ns 2.0V 305360000.0ns 2.0V 305400000.0ns 2.0V 305880000.0ns 2.0V 305920000.0ns 2.0V 306640000.0ns 2.0V 306680000.0ns 0V 307160000.0ns 0V 307200000.0ns 2.0V 307920000.0ns 2.0V 307960000.0ns 2.0V 308440000.0ns 2.0V 308480000.0ns 2.0V 309200000.0ns 2.0V 309240000.0ns 2.0V 309720000.0ns 2.0V 309760000.0ns 2.0V 310480000.0ns 2.0V 310520000.0ns 0V 311000000.0ns 0V 311040000.0ns 2.0V 311760000.0ns 2.0V 311800000.0ns 2.0V 312280000.0ns 2.0V 312320000.0ns 2.0V 313040000.0ns 2.0V 313080000.0ns 2.0V 313560000.0ns 2.0V 313600000.0ns 2.0V 314320000.0ns 2.0V 314360000.0ns 0V 314840000.0ns 0V 314880000.0ns 2.0V 315600000.0ns 2.0V 315640000.0ns 2.0V 316120000.0ns 2.0V 316160000.0ns 2.0V 316880000.0ns 2.0V 316920000.0ns 2.0V 317400000.0ns 2.0V 317440000.0ns 2.0V 318160000.0ns 2.0V 318200000.0ns 0V 318680000.0ns 0V 318720000.0ns 2.0V 319440000.0ns 2.0V 319480000.0ns 2.0V 319960000.0ns 2.0V 320000000.0ns 2.0V 320720000.0ns 2.0V 320760000.0ns 2.0V 321240000.0ns 2.0V 321280000.0ns 2.0V 322000000.0ns 2.0V 322040000.0ns 0V 322520000.0ns 0V 322560000.0ns 2.0V 323280000.0ns 2.0V 323320000.0ns 2.0V 323800000.0ns 2.0V 323840000.0ns 2.0V 324560000.0ns 2.0V 324600000.0ns 2.0V 325080000.0ns 2.0V 325120000.0ns 2.0V 325840000.0ns 2.0V 325880000.0ns 0V 326360000.0ns 0V 326400000.0ns 2.0V 327120000.0ns 2.0V 327160000.0ns 2.0V 327640000.0ns 2.0V 327680000.0ns 2.0V 328400000.0ns 2.0V 328440000.0ns 2.0V 328920000.0ns 2.0V 328960000.0ns 2.0V 329680000.0ns 2.0V 329720000.0ns 0V 330200000.0ns 0V 330240000.0ns 2.0V 330960000.0ns 2.0V 331000000.0ns 2.0V 331480000.0ns 2.0V 331520000.0ns 2.0V 332240000.0ns 2.0V 332280000.0ns 2.0V 332760000.0ns 2.0V 332800000.0ns 2.0V 333520000.0ns 2.0V 333560000.0ns 0V 334040000.0ns 0V 334080000.0ns 2.0V 334800000.0ns 2.0V 334840000.0ns 2.0V 335320000.0ns 2.0V 335360000.0ns 2.0V 336080000.0ns 2.0V 336120000.0ns 2.0V 336600000.0ns 2.0V 336640000.0ns 2.0V 337360000.0ns 2.0V 337400000.0ns 0V 337880000.0ns 0V 337920000.0ns 2.0V 338640000.0ns 2.0V 338680000.0ns 2.0V 339160000.0ns 2.0V 339200000.0ns 2.0V 339920000.0ns 2.0V 339960000.0ns 2.0V 340440000.0ns 2.0V 340480000.0ns 2.0V 341200000.0ns 2.0V 341240000.0ns 0V 341720000.0ns 0V 341760000.0ns 2.0V 342480000.0ns 2.0V 342520000.0ns 2.0V 343000000.0ns 2.0V 343040000.0ns 2.0V 343760000.0ns 2.0V 343800000.0ns 2.0V 344280000.0ns 2.0V 344320000.0ns 2.0V 345040000.0ns 2.0V 345080000.0ns 0V 345560000.0ns 0V 345600000.0ns 2.0V 346320000.0ns 2.0V 346360000.0ns 2.0V 346840000.0ns 2.0V 346880000.0ns 2.0V 347600000.0ns 2.0V 347640000.0ns 2.0V 348120000.0ns 2.0V 348160000.0ns 2.0V 348880000.0ns 2.0V 348920000.0ns 0V 349400000.0ns 0V 349440000.0ns 2.0V 350160000.0ns 2.0V 350200000.0ns 2.0V 350680000.0ns 2.0V 350720000.0ns 2.0V 351440000.0ns 2.0V 351480000.0ns 2.0V 351960000.0ns 2.0V 352000000.0ns 2.0V 352720000.0ns 2.0V 352760000.0ns 0V 353240000.0ns 0V 353280000.0ns 2.0V 354000000.0ns 2.0V 354040000.0ns 2.0V 354520000.0ns 2.0V 354560000.0ns 2.0V 355280000.0ns 2.0V 355320000.0ns 2.0V 355800000.0ns 2.0V 355840000.0ns 2.0V 356560000.0ns 2.0V 356600000.0ns 0V 357080000.0ns 0V 357120000.0ns 2.0V 357840000.0ns 2.0V 357880000.0ns 2.0V 358360000.0ns 2.0V 358400000.0ns 2.0V 359120000.0ns 2.0V 359160000.0ns 2.0V 359640000.0ns 2.0V 359680000.0ns 2.0V 360400000.0ns 2.0V 360440000.0ns 0V 360920000.0ns 0V 360960000.0ns 2.0V 361680000.0ns 2.0V 361720000.0ns 2.0V 362200000.0ns 2.0V 362240000.0ns 2.0V 362960000.0ns 2.0V 363000000.0ns 2.0V 363480000.0ns 2.0V 363520000.0ns 2.0V 364240000.0ns 2.0V 364280000.0ns 0V 364760000.0ns 0V 364800000.0ns 2.0V 365520000.0ns 2.0V 365560000.0ns 2.0V 366040000.0ns 2.0V 366080000.0ns 2.0V 366800000.0ns 2.0V 366840000.0ns 2.0V 367320000.0ns 2.0V 367360000.0ns 2.0V 368080000.0ns 2.0V 368120000.0ns 0V 368600000.0ns 0V 368640000.0ns 2.0V 369360000.0ns 2.0V 369400000.0ns 2.0V 369880000.0ns 2.0V 369920000.0ns 2.0V 370640000.0ns 2.0V 370680000.0ns 2.0V 371160000.0ns 2.0V 371200000.0ns 2.0V 371920000.0ns 2.0V 371960000.0ns 0V 372440000.0ns 0V 372480000.0ns 2.0V 373200000.0ns 2.0V 373240000.0ns 2.0V 373720000.0ns 2.0V 373760000.0ns 2.0V 374480000.0ns 2.0V 374520000.0ns 2.0V 375000000.0ns 2.0V 375040000.0ns 2.0V 375760000.0ns 2.0V 375800000.0ns 0V 376280000.0ns 0V 376320000.0ns 2.0V 377040000.0ns 2.0V 377080000.0ns 2.0V 377560000.0ns 2.0V 377600000.0ns 2.0V 378320000.0ns 2.0V 378360000.0ns 2.0V 378840000.0ns 2.0V 378880000.0ns 2.0V 379600000.0ns 2.0V 379640000.0ns 0V 380120000.0ns 0V 380160000.0ns 2.0V 380880000.0ns 2.0V 380920000.0ns 2.0V 381400000.0ns 2.0V 381440000.0ns 2.0V 382160000.0ns 2.0V 382200000.0ns 2.0V 382680000.0ns 2.0V 382720000.0ns 2.0V 383440000.0ns 2.0V 383480000.0ns 0V 383960000.0ns 0V 384000000.0ns 2.0V 384720000.0ns 2.0V 384760000.0ns 2.0V 385240000.0ns 2.0V 385280000.0ns 2.0V 386000000.0ns 2.0V 386040000.0ns 2.0V 386520000.0ns 2.0V 386560000.0ns 2.0V 387280000.0ns 2.0V 387320000.0ns 0V 387800000.0ns 0V 387840000.0ns 2.0V 388560000.0ns 2.0V 388600000.0ns 2.0V 389080000.0ns 2.0V 389120000.0ns 2.0V 389840000.0ns 2.0V 389880000.0ns 2.0V 390360000.0ns 2.0V 390400000.0ns 2.0V 391120000.0ns 2.0V 391160000.0ns 0V)
Vtarget_0 target_0 0 PWL(0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0.27862048149108887V 8400000.0ns 0.27862048149108887V 8440000.0ns 0.27862048149108887V 8920000.0ns 0.27862048149108887V 8960000.0ns 0.27862048149108887V 9680000.0ns 0.27862048149108887V 9720000.0ns 0.27862048149108887V 10200000.0ns 0.27862048149108887V 10240000.0ns 0.27862048149108887V 10960000.0ns 0.27862048149108887V 11000000.0ns 0V 11480000.0ns 0V 11520000.0ns 0.29986271262168884V 12240000.0ns 0.29986271262168884V 12280000.0ns 0.29986271262168884V 12760000.0ns 0.29986271262168884V 12800000.0ns 0.29986271262168884V 13520000.0ns 0.29986271262168884V 13560000.0ns 0.29986271262168884V 14040000.0ns 0.29986271262168884V 14080000.0ns 0.29986271262168884V 14800000.0ns 0.29986271262168884V 14840000.0ns 0V 15320000.0ns 0V 15360000.0ns 0.15744949877262115V 16080000.0ns 0.15744949877262115V 16120000.0ns 0.15744949877262115V 16600000.0ns 0.15744949877262115V 16640000.0ns 0.15744949877262115V 17360000.0ns 0.15744949877262115V 17400000.0ns 0.15744949877262115V 17880000.0ns 0.15744949877262115V 17920000.0ns 0.15744949877262115V 18640000.0ns 0.15744949877262115V 18680000.0ns 0V 19160000.0ns 0V 19200000.0ns 0.10012375563383102V 19920000.0ns 0.10012375563383102V 19960000.0ns 0.10012375563383102V 20440000.0ns 0.10012375563383102V 20480000.0ns 0.10012375563383102V 21200000.0ns 0.10012375563383102V 21240000.0ns 0.10012375563383102V 21720000.0ns 0.10012375563383102V 21760000.0ns 0.10012375563383102V 22480000.0ns 0.10012375563383102V 22520000.0ns 0V 23000000.0ns 0V 23040000.0ns 0.29320797324180603V 23760000.0ns 0.29320797324180603V 23800000.0ns 0.29320797324180603V 24280000.0ns 0.29320797324180603V 24320000.0ns 0.29320797324180603V 25040000.0ns 0.29320797324180603V 25080000.0ns 0.29320797324180603V 25560000.0ns 0.29320797324180603V 25600000.0ns 0.29320797324180603V 26320000.0ns 0.29320797324180603V 26360000.0ns 0V 26840000.0ns 0V 26880000.0ns 0.23135295510292053V 27600000.0ns 0.23135295510292053V 27640000.0ns 0.23135295510292053V 28120000.0ns 0.23135295510292053V 28160000.0ns 0.23135295510292053V 28880000.0ns 0.23135295510292053V 28920000.0ns 0.23135295510292053V 29400000.0ns 0.23135295510292053V 29440000.0ns 0.23135295510292053V 30160000.0ns 0.23135295510292053V 30200000.0ns 0V 30680000.0ns 0V 30720000.0ns 0.2570348083972931V 31440000.0ns 0.2570348083972931V 31480000.0ns 0.2570348083972931V 31960000.0ns 0.2570348083972931V 32000000.0ns 0.2570348083972931V 32720000.0ns 0.2570348083972931V 32760000.0ns 0.2570348083972931V 33240000.0ns 0.2570348083972931V 33280000.0ns 0.2570348083972931V 34000000.0ns 0.2570348083972931V 34040000.0ns 0V 34520000.0ns 0V 34560000.0ns 0.157086580991745V 35280000.0ns 0.157086580991745V 35320000.0ns 0.157086580991745V 35800000.0ns 0.157086580991745V 35840000.0ns 0.157086580991745V 36560000.0ns 0.157086580991745V 36600000.0ns 0.157086580991745V 37080000.0ns 0.157086580991745V 37120000.0ns 0.157086580991745V 37840000.0ns 0.157086580991745V 37880000.0ns 0V 38360000.0ns 0V 38400000.0ns 0.23427122831344604V 39120000.0ns 0.23427122831344604V 39160000.0ns 0.23427122831344604V 39640000.0ns 0.23427122831344604V 39680000.0ns 0.23427122831344604V 40400000.0ns 0.23427122831344604V 40440000.0ns 0.23427122831344604V 40920000.0ns 0.23427122831344604V 40960000.0ns 0.23427122831344604V 41680000.0ns 0.23427122831344604V 41720000.0ns 0V 42200000.0ns 0V 42240000.0ns 0.26756608486175537V 42960000.0ns 0.26756608486175537V 43000000.0ns 0.26756608486175537V 43480000.0ns 0.26756608486175537V 43520000.0ns 0.26756608486175537V 44240000.0ns 0.26756608486175537V 44280000.0ns 0.26756608486175537V 44760000.0ns 0.26756608486175537V 44800000.0ns 0.26756608486175537V 45520000.0ns 0.26756608486175537V 45560000.0ns 0V 46040000.0ns 0V 46080000.0ns 0.2859998047351837V 46800000.0ns 0.2859998047351837V 46840000.0ns 0.2859998047351837V 47320000.0ns 0.2859998047351837V 47360000.0ns 0.2859998047351837V 48080000.0ns 0.2859998047351837V 48120000.0ns 0.2859998047351837V 48600000.0ns 0.2859998047351837V 48640000.0ns 0.2859998047351837V 49360000.0ns 0.2859998047351837V 49400000.0ns 0V 49880000.0ns 0V 49920000.0ns 0.18126188218593597V 50640000.0ns 0.18126188218593597V 50680000.0ns 0.18126188218593597V 51160000.0ns 0.18126188218593597V 51200000.0ns 0.18126188218593597V 51920000.0ns 0.18126188218593597V 51960000.0ns 0.18126188218593597V 52440000.0ns 0.18126188218593597V 52480000.0ns 0.18126188218593597V 53200000.0ns 0.18126188218593597V 53240000.0ns 0V 53720000.0ns 0V 53760000.0ns 0.2565646469593048V 54480000.0ns 0.2565646469593048V 54520000.0ns 0.2565646469593048V 55000000.0ns 0.2565646469593048V 55040000.0ns 0.2565646469593048V 55760000.0ns 0.2565646469593048V 55800000.0ns 0.2565646469593048V 56280000.0ns 0.2565646469593048V 56320000.0ns 0.2565646469593048V 57040000.0ns 0.2565646469593048V 57080000.0ns 0V 57560000.0ns 0V 57600000.0ns 0.2732909917831421V 58320000.0ns 0.2732909917831421V 58360000.0ns 0.2732909917831421V 58840000.0ns 0.2732909917831421V 58880000.0ns 0.2732909917831421V 59600000.0ns 0.2732909917831421V 59640000.0ns 0.2732909917831421V 60120000.0ns 0.2732909917831421V 60160000.0ns 0.2732909917831421V 60880000.0ns 0.2732909917831421V 60920000.0ns 0V 61400000.0ns 0V 61440000.0ns 0.17634646594524384V 62160000.0ns 0.17634646594524384V 62200000.0ns 0.17634646594524384V 62680000.0ns 0.17634646594524384V 62720000.0ns 0.17634646594524384V 63440000.0ns 0.17634646594524384V 63480000.0ns 0.17634646594524384V 63960000.0ns 0.17634646594524384V 64000000.0ns 0.17634646594524384V 64720000.0ns 0.17634646594524384V 64760000.0ns 0V 65240000.0ns 0V 65280000.0ns 0.12059792876243591V 66000000.0ns 0.12059792876243591V 66040000.0ns 0.12059792876243591V 66520000.0ns 0.12059792876243591V 66560000.0ns 0.12059792876243591V 67280000.0ns 0.12059792876243591V 67320000.0ns 0.12059792876243591V 67800000.0ns 0.12059792876243591V 67840000.0ns 0.12059792876243591V 68560000.0ns 0.12059792876243591V 68600000.0ns 0V 69080000.0ns 0V 69120000.0ns 0.11544250696897507V 69840000.0ns 0.11544250696897507V 69880000.0ns 0.11544250696897507V 70360000.0ns 0.11544250696897507V 70400000.0ns 0.11544250696897507V 71120000.0ns 0.11544250696897507V 71160000.0ns 0.11544250696897507V 71640000.0ns 0.11544250696897507V 71680000.0ns 0.11544250696897507V 72400000.0ns 0.11544250696897507V 72440000.0ns 0V 72920000.0ns 0V 72960000.0ns 0.14201870560646057V 73680000.0ns 0.14201870560646057V 73720000.0ns 0.14201870560646057V 74200000.0ns 0.14201870560646057V 74240000.0ns 0.14201870560646057V 74960000.0ns 0.14201870560646057V 75000000.0ns 0.14201870560646057V 75480000.0ns 0.14201870560646057V 75520000.0ns 0.14201870560646057V 76240000.0ns 0.14201870560646057V 76280000.0ns 0V 76760000.0ns 0V 76800000.0ns 0.28229114413261414V 77520000.0ns 0.28229114413261414V 77560000.0ns 0.28229114413261414V 78040000.0ns 0.28229114413261414V 78080000.0ns 0.28229114413261414V 78800000.0ns 0.28229114413261414V 78840000.0ns 0.28229114413261414V 79320000.0ns 0.28229114413261414V 79360000.0ns 0.28229114413261414V 80080000.0ns 0.28229114413261414V 80120000.0ns 0V 80600000.0ns 0V 80640000.0ns 0.2995724678039551V 81360000.0ns 0.2995724678039551V 81400000.0ns 0.2995724678039551V 81880000.0ns 0.2995724678039551V 81920000.0ns 0.2995724678039551V 82640000.0ns 0.2995724678039551V 82680000.0ns 0.2995724678039551V 83160000.0ns 0.2995724678039551V 83200000.0ns 0.2995724678039551V 83920000.0ns 0.2995724678039551V 83960000.0ns 0V 84440000.0ns 0V 84480000.0ns 0.2989230155944824V 85200000.0ns 0.2989230155944824V 85240000.0ns 0.2989230155944824V 85720000.0ns 0.2989230155944824V 85760000.0ns 0.2989230155944824V 86480000.0ns 0.2989230155944824V 86520000.0ns 0.2989230155944824V 87000000.0ns 0.2989230155944824V 87040000.0ns 0.2989230155944824V 87760000.0ns 0.2989230155944824V 87800000.0ns 0V 88280000.0ns 0V 88320000.0ns 0.2903580665588379V 89040000.0ns 0.2903580665588379V 89080000.0ns 0.2903580665588379V 89560000.0ns 0.2903580665588379V 89600000.0ns 0.2903580665588379V 90320000.0ns 0.2903580665588379V 90360000.0ns 0.2903580665588379V 90840000.0ns 0.2903580665588379V 90880000.0ns 0.2903580665588379V 91600000.0ns 0.2903580665588379V 91640000.0ns 0V 92120000.0ns 0V 92160000.0ns 0.24801762402057648V 92880000.0ns 0.24801762402057648V 92920000.0ns 0.24801762402057648V 93400000.0ns 0.24801762402057648V 93440000.0ns 0.24801762402057648V 94160000.0ns 0.24801762402057648V 94200000.0ns 0.24801762402057648V 94680000.0ns 0.24801762402057648V 94720000.0ns 0.24801762402057648V 95440000.0ns 0.24801762402057648V 95480000.0ns 0V 95960000.0ns 0V 96000000.0ns 0.26778000593185425V 96720000.0ns 0.26778000593185425V 96760000.0ns 0.26778000593185425V 97240000.0ns 0.26778000593185425V 97280000.0ns 0.26778000593185425V 98000000.0ns 0.26778000593185425V 98040000.0ns 0.26778000593185425V 98520000.0ns 0.26778000593185425V 98560000.0ns 0.26778000593185425V 99280000.0ns 0.26778000593185425V 99320000.0ns 0V 99800000.0ns 0V 99840000.0ns 0.12881134450435638V 100560000.0ns 0.12881134450435638V 100600000.0ns 0.12881134450435638V 101080000.0ns 0.12881134450435638V 101120000.0ns 0.12881134450435638V 101840000.0ns 0.12881134450435638V 101880000.0ns 0.12881134450435638V 102360000.0ns 0.12881134450435638V 102400000.0ns 0.12881134450435638V 103120000.0ns 0.12881134450435638V 103160000.0ns 0V 103640000.0ns 0V 103680000.0ns 0.20720621943473816V 104400000.0ns 0.20720621943473816V 104440000.0ns 0.20720621943473816V 104920000.0ns 0.20720621943473816V 104960000.0ns 0.20720621943473816V 105680000.0ns 0.20720621943473816V 105720000.0ns 0.20720621943473816V 106200000.0ns 0.20720621943473816V 106240000.0ns 0.20720621943473816V 106960000.0ns 0.20720621943473816V 107000000.0ns 0V 107480000.0ns 0V 107520000.0ns 0.22566945850849152V 108240000.0ns 0.22566945850849152V 108280000.0ns 0.22566945850849152V 108760000.0ns 0.22566945850849152V 108800000.0ns 0.22566945850849152V 109520000.0ns 0.22566945850849152V 109560000.0ns 0.22566945850849152V 110040000.0ns 0.22566945850849152V 110080000.0ns 0.22566945850849152V 110800000.0ns 0.22566945850849152V 110840000.0ns 0V 111320000.0ns 0V 111360000.0ns 0.24488961696624756V 112080000.0ns 0.24488961696624756V 112120000.0ns 0.24488961696624756V 112600000.0ns 0.24488961696624756V 112640000.0ns 0.24488961696624756V 113360000.0ns 0.24488961696624756V 113400000.0ns 0.24488961696624756V 113880000.0ns 0.24488961696624756V 113920000.0ns 0.24488961696624756V 114640000.0ns 0.24488961696624756V 114680000.0ns 0V 115160000.0ns 0V 115200000.0ns 0.2678714394569397V 115920000.0ns 0.2678714394569397V 115960000.0ns 0.2678714394569397V 116440000.0ns 0.2678714394569397V 116480000.0ns 0.2678714394569397V 117200000.0ns 0.2678714394569397V 117240000.0ns 0.2678714394569397V 117720000.0ns 0.2678714394569397V 117760000.0ns 0.2678714394569397V 118480000.0ns 0.2678714394569397V 118520000.0ns 0V 119000000.0ns 0V 119040000.0ns 0.19972366094589233V 119760000.0ns 0.19972366094589233V 119800000.0ns 0.19972366094589233V 120280000.0ns 0.19972366094589233V 120320000.0ns 0.19972366094589233V 121040000.0ns 0.19972366094589233V 121080000.0ns 0.19972366094589233V 121560000.0ns 0.19972366094589233V 121600000.0ns 0.19972366094589233V 122320000.0ns 0.19972366094589233V 122360000.0ns 0V 122840000.0ns 0V 122880000.0ns 0.2868887782096863V 123600000.0ns 0.2868887782096863V 123640000.0ns 0.2868887782096863V 124120000.0ns 0.2868887782096863V 124160000.0ns 0.2868887782096863V 124880000.0ns 0.2868887782096863V 124920000.0ns 0.2868887782096863V 125400000.0ns 0.2868887782096863V 125440000.0ns 0.2868887782096863V 126160000.0ns 0.2868887782096863V 126200000.0ns 0V 126680000.0ns 0V 126720000.0ns 0.10920276492834091V 127440000.0ns 0.10920276492834091V 127480000.0ns 0.10920276492834091V 127960000.0ns 0.10920276492834091V 128000000.0ns 0.10920276492834091V 128720000.0ns 0.10920276492834091V 128760000.0ns 0.10920276492834091V 129240000.0ns 0.10920276492834091V 129280000.0ns 0.10920276492834091V 130000000.0ns 0.10920276492834091V 130040000.0ns 0V 130520000.0ns 0V 130560000.0ns 0.21748633682727814V 131280000.0ns 0.21748633682727814V 131320000.0ns 0.21748633682727814V 131800000.0ns 0.21748633682727814V 131840000.0ns 0.21748633682727814V 132560000.0ns 0.21748633682727814V 132600000.0ns 0.21748633682727814V 133080000.0ns 0.21748633682727814V 133120000.0ns 0.21748633682727814V 133840000.0ns 0.21748633682727814V 133880000.0ns 0V 134360000.0ns 0V 134400000.0ns 0.25955140590667725V 135120000.0ns 0.25955140590667725V 135160000.0ns 0.25955140590667725V 135640000.0ns 0.25955140590667725V 135680000.0ns 0.25955140590667725V 136400000.0ns 0.25955140590667725V 136440000.0ns 0.25955140590667725V 136920000.0ns 0.25955140590667725V 136960000.0ns 0.25955140590667725V 137680000.0ns 0.25955140590667725V 137720000.0ns 0V 138200000.0ns 0V 138240000.0ns 0.2493583709001541V 138960000.0ns 0.2493583709001541V 139000000.0ns 0.2493583709001541V 139480000.0ns 0.2493583709001541V 139520000.0ns 0.2493583709001541V 140240000.0ns 0.2493583709001541V 140280000.0ns 0.2493583709001541V 140760000.0ns 0.2493583709001541V 140800000.0ns 0.2493583709001541V 141520000.0ns 0.2493583709001541V 141560000.0ns 0V 142040000.0ns 0V 142080000.0ns 0.2994815707206726V 142800000.0ns 0.2994815707206726V 142840000.0ns 0.2994815707206726V 143320000.0ns 0.2994815707206726V 143360000.0ns 0.2994815707206726V 144080000.0ns 0.2994815707206726V 144120000.0ns 0.2994815707206726V 144600000.0ns 0.2994815707206726V 144640000.0ns 0.2994815707206726V 145360000.0ns 0.2994815707206726V 145400000.0ns 0V 145880000.0ns 0V 145920000.0ns 0.11542080342769623V 146640000.0ns 0.11542080342769623V 146680000.0ns 0.11542080342769623V 147160000.0ns 0.11542080342769623V 147200000.0ns 0.11542080342769623V 147920000.0ns 0.11542080342769623V 147960000.0ns 0.11542080342769623V 148440000.0ns 0.11542080342769623V 148480000.0ns 0.11542080342769623V 149200000.0ns 0.11542080342769623V 149240000.0ns 0V 149720000.0ns 0V 149760000.0ns 0.299551397562027V 150480000.0ns 0.299551397562027V 150520000.0ns 0.299551397562027V 151000000.0ns 0.299551397562027V 151040000.0ns 0.299551397562027V 151760000.0ns 0.299551397562027V 151800000.0ns 0.299551397562027V 152280000.0ns 0.299551397562027V 152320000.0ns 0.299551397562027V 153040000.0ns 0.299551397562027V 153080000.0ns 0V 153560000.0ns 0V 153600000.0ns 0.1503254473209381V 154320000.0ns 0.1503254473209381V 154360000.0ns 0.1503254473209381V 154840000.0ns 0.1503254473209381V 154880000.0ns 0.1503254473209381V 155600000.0ns 0.1503254473209381V 155640000.0ns 0.1503254473209381V 156120000.0ns 0.1503254473209381V 156160000.0ns 0.1503254473209381V 156880000.0ns 0.1503254473209381V 156920000.0ns 0V 157400000.0ns 0V 157440000.0ns 0.29132726788520813V 158160000.0ns 0.29132726788520813V 158200000.0ns 0.29132726788520813V 158680000.0ns 0.29132726788520813V 158720000.0ns 0.29132726788520813V 159440000.0ns 0.29132726788520813V 159480000.0ns 0.29132726788520813V 159960000.0ns 0.29132726788520813V 160000000.0ns 0.29132726788520813V 160720000.0ns 0.29132726788520813V 160760000.0ns 0V 161240000.0ns 0V 161280000.0ns 0.2605951428413391V 162000000.0ns 0.2605951428413391V 162040000.0ns 0.2605951428413391V 162520000.0ns 0.2605951428413391V 162560000.0ns 0.2605951428413391V 163280000.0ns 0.2605951428413391V 163320000.0ns 0.2605951428413391V 163800000.0ns 0.2605951428413391V 163840000.0ns 0.2605951428413391V 164560000.0ns 0.2605951428413391V 164600000.0ns 0V 165080000.0ns 0V 165120000.0ns 0.29995816946029663V 165840000.0ns 0.29995816946029663V 165880000.0ns 0.29995816946029663V 166360000.0ns 0.29995816946029663V 166400000.0ns 0.29995816946029663V 167120000.0ns 0.29995816946029663V 167160000.0ns 0.29995816946029663V 167640000.0ns 0.29995816946029663V 167680000.0ns 0.29995816946029663V 168400000.0ns 0.29995816946029663V 168440000.0ns 0V 168920000.0ns 0V 168960000.0ns 0.2621794641017914V 169680000.0ns 0.2621794641017914V 169720000.0ns 0.2621794641017914V 170200000.0ns 0.2621794641017914V 170240000.0ns 0.2621794641017914V 170960000.0ns 0.2621794641017914V 171000000.0ns 0.2621794641017914V 171480000.0ns 0.2621794641017914V 171520000.0ns 0.2621794641017914V 172240000.0ns 0.2621794641017914V 172280000.0ns 0V 172760000.0ns 0V 172800000.0ns 0.2382839322090149V 173520000.0ns 0.2382839322090149V 173560000.0ns 0.2382839322090149V 174040000.0ns 0.2382839322090149V 174080000.0ns 0.2382839322090149V 174800000.0ns 0.2382839322090149V 174840000.0ns 0.2382839322090149V 175320000.0ns 0.2382839322090149V 175360000.0ns 0.2382839322090149V 176080000.0ns 0.2382839322090149V 176120000.0ns 0V 176600000.0ns 0V 176640000.0ns 0.1269591748714447V 177360000.0ns 0.1269591748714447V 177400000.0ns 0.1269591748714447V 177880000.0ns 0.1269591748714447V 177920000.0ns 0.1269591748714447V 178640000.0ns 0.1269591748714447V 178680000.0ns 0.1269591748714447V 179160000.0ns 0.1269591748714447V 179200000.0ns 0.1269591748714447V 179920000.0ns 0.1269591748714447V 179960000.0ns 0V 180440000.0ns 0V 180480000.0ns 0.10124511271715164V 181200000.0ns 0.10124511271715164V 181240000.0ns 0.10124511271715164V 181720000.0ns 0.10124511271715164V 181760000.0ns 0.10124511271715164V 182480000.0ns 0.10124511271715164V 182520000.0ns 0.10124511271715164V 183000000.0ns 0.10124511271715164V 183040000.0ns 0.10124511271715164V 183760000.0ns 0.10124511271715164V 183800000.0ns 0V 184280000.0ns 0V 184320000.0ns 0.22850382328033447V 185040000.0ns 0.22850382328033447V 185080000.0ns 0.22850382328033447V 185560000.0ns 0.22850382328033447V 185600000.0ns 0.22850382328033447V 186320000.0ns 0.22850382328033447V 186360000.0ns 0.22850382328033447V 186840000.0ns 0.22850382328033447V 186880000.0ns 0.22850382328033447V 187600000.0ns 0.22850382328033447V 187640000.0ns 0V 188120000.0ns 0V 188160000.0ns 0.10704908519983292V 188880000.0ns 0.10704908519983292V 188920000.0ns 0.10704908519983292V 189400000.0ns 0.10704908519983292V 189440000.0ns 0.10704908519983292V 190160000.0ns 0.10704908519983292V 190200000.0ns 0.10704908519983292V 190680000.0ns 0.10704908519983292V 190720000.0ns 0.10704908519983292V 191440000.0ns 0.10704908519983292V 191480000.0ns 0V 191960000.0ns 0V 192000000.0ns 0.22501061856746674V 192720000.0ns 0.22501061856746674V 192760000.0ns 0.22501061856746674V 193240000.0ns 0.22501061856746674V 193280000.0ns 0.22501061856746674V 194000000.0ns 0.22501061856746674V 194040000.0ns 0.22501061856746674V 194520000.0ns 0.22501061856746674V 194560000.0ns 0.22501061856746674V 195280000.0ns 0.22501061856746674V 195320000.0ns 0V 195800000.0ns 0V 195840000.0ns 0.2122419774532318V 196560000.0ns 0.2122419774532318V 196600000.0ns 0.2122419774532318V 197080000.0ns 0.2122419774532318V 197120000.0ns 0.2122419774532318V 197840000.0ns 0.2122419774532318V 197880000.0ns 0.2122419774532318V 198360000.0ns 0.2122419774532318V 198400000.0ns 0.2122419774532318V 199120000.0ns 0.2122419774532318V 199160000.0ns 0V 199640000.0ns 0V 199680000.0ns 0.29918158054351807V 200400000.0ns 0.29918158054351807V 200440000.0ns 0.29918158054351807V 200920000.0ns 0.29918158054351807V 200960000.0ns 0.29918158054351807V 201680000.0ns 0.29918158054351807V 201720000.0ns 0.29918158054351807V 202200000.0ns 0.29918158054351807V 202240000.0ns 0.29918158054351807V 202960000.0ns 0.29918158054351807V 203000000.0ns 0V 203480000.0ns 0V 203520000.0ns 0.10419157892465591V 204240000.0ns 0.10419157892465591V 204280000.0ns 0.10419157892465591V 204760000.0ns 0.10419157892465591V 204800000.0ns 0.10419157892465591V 205520000.0ns 0.10419157892465591V 205560000.0ns 0.10419157892465591V 206040000.0ns 0.10419157892465591V 206080000.0ns 0.10419157892465591V 206800000.0ns 0.10419157892465591V 206840000.0ns 0V 207320000.0ns 0V 207360000.0ns 0.1528206467628479V 208080000.0ns 0.1528206467628479V 208120000.0ns 0.1528206467628479V 208600000.0ns 0.1528206467628479V 208640000.0ns 0.1528206467628479V 209360000.0ns 0.1528206467628479V 209400000.0ns 0.1528206467628479V 209880000.0ns 0.1528206467628479V 209920000.0ns 0.1528206467628479V 210640000.0ns 0.1528206467628479V 210680000.0ns 0V 211160000.0ns 0V 211200000.0ns 0.2971463203430176V 211920000.0ns 0.2971463203430176V 211960000.0ns 0.2971463203430176V 212440000.0ns 0.2971463203430176V 212480000.0ns 0.2971463203430176V 213200000.0ns 0.2971463203430176V 213240000.0ns 0.2971463203430176V 213720000.0ns 0.2971463203430176V 213760000.0ns 0.2971463203430176V 214480000.0ns 0.2971463203430176V 214520000.0ns 0V 215000000.0ns 0V 215040000.0ns 0.17168807983398438V 215760000.0ns 0.17168807983398438V 215800000.0ns 0.17168807983398438V 216280000.0ns 0.17168807983398438V 216320000.0ns 0.17168807983398438V 217040000.0ns 0.17168807983398438V 217080000.0ns 0.17168807983398438V 217560000.0ns 0.17168807983398438V 217600000.0ns 0.17168807983398438V 218320000.0ns 0.17168807983398438V 218360000.0ns 0V 218840000.0ns 0V 218880000.0ns 0.2648089826107025V 219600000.0ns 0.2648089826107025V 219640000.0ns 0.2648089826107025V 220120000.0ns 0.2648089826107025V 220160000.0ns 0.2648089826107025V 220880000.0ns 0.2648089826107025V 220920000.0ns 0.2648089826107025V 221400000.0ns 0.2648089826107025V 221440000.0ns 0.2648089826107025V 222160000.0ns 0.2648089826107025V 222200000.0ns 0V 222680000.0ns 0V 222720000.0ns 0.2902770936489105V 223440000.0ns 0.2902770936489105V 223480000.0ns 0.2902770936489105V 223960000.0ns 0.2902770936489105V 224000000.0ns 0.2902770936489105V 224720000.0ns 0.2902770936489105V 224760000.0ns 0.2902770936489105V 225240000.0ns 0.2902770936489105V 225280000.0ns 0.2902770936489105V 226000000.0ns 0.2902770936489105V 226040000.0ns 0V 226520000.0ns 0V 226560000.0ns 0.19853074848651886V 227280000.0ns 0.19853074848651886V 227320000.0ns 0.19853074848651886V 227800000.0ns 0.19853074848651886V 227840000.0ns 0.19853074848651886V 228560000.0ns 0.19853074848651886V 228600000.0ns 0.19853074848651886V 229080000.0ns 0.19853074848651886V 229120000.0ns 0.19853074848651886V 229840000.0ns 0.19853074848651886V 229880000.0ns 0V 230360000.0ns 0V 230400000.0ns 0.21381524205207825V 231120000.0ns 0.21381524205207825V 231160000.0ns 0.21381524205207825V 231640000.0ns 0.21381524205207825V 231680000.0ns 0.21381524205207825V 232400000.0ns 0.21381524205207825V 232440000.0ns 0.21381524205207825V 232920000.0ns 0.21381524205207825V 232960000.0ns 0.21381524205207825V 233680000.0ns 0.21381524205207825V 233720000.0ns 0V 234200000.0ns 0V 234240000.0ns 0.26878055930137634V 234960000.0ns 0.26878055930137634V 235000000.0ns 0.26878055930137634V 235480000.0ns 0.26878055930137634V 235520000.0ns 0.26878055930137634V 236240000.0ns 0.26878055930137634V 236280000.0ns 0.26878055930137634V 236760000.0ns 0.26878055930137634V 236800000.0ns 0.26878055930137634V 237520000.0ns 0.26878055930137634V 237560000.0ns 0V 238040000.0ns 0V 238080000.0ns 0.20533791184425354V 238800000.0ns 0.20533791184425354V 238840000.0ns 0.20533791184425354V 239320000.0ns 0.20533791184425354V 239360000.0ns 0.20533791184425354V 240080000.0ns 0.20533791184425354V 240120000.0ns 0.20533791184425354V 240600000.0ns 0.20533791184425354V 240640000.0ns 0.20533791184425354V 241360000.0ns 0.20533791184425354V 241400000.0ns 0V 241880000.0ns 0V 241920000.0ns 0.23522275686264038V 242640000.0ns 0.23522275686264038V 242680000.0ns 0.23522275686264038V 243160000.0ns 0.23522275686264038V 243200000.0ns 0.23522275686264038V 243920000.0ns 0.23522275686264038V 243960000.0ns 0.23522275686264038V 244440000.0ns 0.23522275686264038V 244480000.0ns 0.23522275686264038V 245200000.0ns 0.23522275686264038V 245240000.0ns 0V 245720000.0ns 0V 245760000.0ns 0.29486843943595886V 246480000.0ns 0.29486843943595886V 246520000.0ns 0.29486843943595886V 247000000.0ns 0.29486843943595886V 247040000.0ns 0.29486843943595886V 247760000.0ns 0.29486843943595886V 247800000.0ns 0.29486843943595886V 248280000.0ns 0.29486843943595886V 248320000.0ns 0.29486843943595886V 249040000.0ns 0.29486843943595886V 249080000.0ns 0V 249560000.0ns 0V 249600000.0ns 0.19978351891040802V 250320000.0ns 0.19978351891040802V 250360000.0ns 0.19978351891040802V 250840000.0ns 0.19978351891040802V 250880000.0ns 0.19978351891040802V 251600000.0ns 0.19978351891040802V 251640000.0ns 0.19978351891040802V 252120000.0ns 0.19978351891040802V 252160000.0ns 0.19978351891040802V 252880000.0ns 0.19978351891040802V 252920000.0ns 0V 253400000.0ns 0V 253440000.0ns 0.174158975481987V 254160000.0ns 0.174158975481987V 254200000.0ns 0.174158975481987V 254680000.0ns 0.174158975481987V 254720000.0ns 0.174158975481987V 255440000.0ns 0.174158975481987V 255480000.0ns 0.174158975481987V 255960000.0ns 0.174158975481987V 256000000.0ns 0.174158975481987V 256720000.0ns 0.174158975481987V 256760000.0ns 0V 257240000.0ns 0V 257280000.0ns 0.18191738426685333V 258000000.0ns 0.18191738426685333V 258040000.0ns 0.18191738426685333V 258520000.0ns 0.18191738426685333V 258560000.0ns 0.18191738426685333V 259280000.0ns 0.18191738426685333V 259320000.0ns 0.18191738426685333V 259800000.0ns 0.18191738426685333V 259840000.0ns 0.18191738426685333V 260560000.0ns 0.18191738426685333V 260600000.0ns 0V 261080000.0ns 0V 261120000.0ns 0.18075774610042572V 261840000.0ns 0.18075774610042572V 261880000.0ns 0.18075774610042572V 262360000.0ns 0.18075774610042572V 262400000.0ns 0.18075774610042572V 263120000.0ns 0.18075774610042572V 263160000.0ns 0.18075774610042572V 263640000.0ns 0.18075774610042572V 263680000.0ns 0.18075774610042572V 264400000.0ns 0.18075774610042572V 264440000.0ns 0V 264920000.0ns 0V 264960000.0ns 0.11365003138780594V 265680000.0ns 0.11365003138780594V 265720000.0ns 0.11365003138780594V 266200000.0ns 0.11365003138780594V 266240000.0ns 0.11365003138780594V 266960000.0ns 0.11365003138780594V 267000000.0ns 0.11365003138780594V 267480000.0ns 0.11365003138780594V 267520000.0ns 0.11365003138780594V 268240000.0ns 0.11365003138780594V 268280000.0ns 0V 268760000.0ns 0V 268800000.0ns 0.18851272761821747V 269520000.0ns 0.18851272761821747V 269560000.0ns 0.18851272761821747V 270040000.0ns 0.18851272761821747V 270080000.0ns 0.18851272761821747V 270800000.0ns 0.18851272761821747V 270840000.0ns 0.18851272761821747V 271320000.0ns 0.18851272761821747V 271360000.0ns 0.18851272761821747V 272080000.0ns 0.18851272761821747V 272120000.0ns 0V 272600000.0ns 0V 272640000.0ns 0.2992361783981323V 273360000.0ns 0.2992361783981323V 273400000.0ns 0.2992361783981323V 273880000.0ns 0.2992361783981323V 273920000.0ns 0.2992361783981323V 274640000.0ns 0.2992361783981323V 274680000.0ns 0.2992361783981323V 275160000.0ns 0.2992361783981323V 275200000.0ns 0.2992361783981323V 275920000.0ns 0.2992361783981323V 275960000.0ns 0V 276440000.0ns 0V 276480000.0ns 0.2109602391719818V 277200000.0ns 0.2109602391719818V 277240000.0ns 0.2109602391719818V 277720000.0ns 0.2109602391719818V 277760000.0ns 0.2109602391719818V 278480000.0ns 0.2109602391719818V 278520000.0ns 0.2109602391719818V 279000000.0ns 0.2109602391719818V 279040000.0ns 0.2109602391719818V 279760000.0ns 0.2109602391719818V 279800000.0ns 0V 280280000.0ns 0V 280320000.0ns 0.2531076669692993V 281040000.0ns 0.2531076669692993V 281080000.0ns 0.2531076669692993V 281560000.0ns 0.2531076669692993V 281600000.0ns 0.2531076669692993V 282320000.0ns 0.2531076669692993V 282360000.0ns 0.2531076669692993V 282840000.0ns 0.2531076669692993V 282880000.0ns 0.2531076669692993V 283600000.0ns 0.2531076669692993V 283640000.0ns 0V 284120000.0ns 0V 284160000.0ns 0.297838032245636V 284880000.0ns 0.297838032245636V 284920000.0ns 0.297838032245636V 285400000.0ns 0.297838032245636V 285440000.0ns 0.297838032245636V 286160000.0ns 0.297838032245636V 286200000.0ns 0.297838032245636V 286680000.0ns 0.297838032245636V 286720000.0ns 0.297838032245636V 287440000.0ns 0.297838032245636V 287480000.0ns 0V 287960000.0ns 0V 288000000.0ns 0.1091398298740387V 288720000.0ns 0.1091398298740387V 288760000.0ns 0.1091398298740387V 289240000.0ns 0.1091398298740387V 289280000.0ns 0.1091398298740387V 290000000.0ns 0.1091398298740387V 290040000.0ns 0.1091398298740387V 290520000.0ns 0.1091398298740387V 290560000.0ns 0.1091398298740387V 291280000.0ns 0.1091398298740387V 291320000.0ns 0V 291800000.0ns 0V 291840000.0ns 0.10169992595911026V 292560000.0ns 0.10169992595911026V 292600000.0ns 0.10169992595911026V 293080000.0ns 0.10169992595911026V 293120000.0ns 0.10169992595911026V 293840000.0ns 0.10169992595911026V 293880000.0ns 0.10169992595911026V 294360000.0ns 0.10169992595911026V 294400000.0ns 0.10169992595911026V 295120000.0ns 0.10169992595911026V 295160000.0ns 0V 295640000.0ns 0V 295680000.0ns 0.12655246257781982V 296400000.0ns 0.12655246257781982V 296440000.0ns 0.12655246257781982V 296920000.0ns 0.12655246257781982V 296960000.0ns 0.12655246257781982V 297680000.0ns 0.12655246257781982V 297720000.0ns 0.12655246257781982V 298200000.0ns 0.12655246257781982V 298240000.0ns 0.12655246257781982V 298960000.0ns 0.12655246257781982V 299000000.0ns 0V 299480000.0ns 0V 299520000.0ns 0.210767462849617V 300240000.0ns 0.210767462849617V 300280000.0ns 0.210767462849617V 300760000.0ns 0.210767462849617V 300800000.0ns 0.210767462849617V 301520000.0ns 0.210767462849617V 301560000.0ns 0.210767462849617V 302040000.0ns 0.210767462849617V 302080000.0ns 0.210767462849617V 302800000.0ns 0.210767462849617V 302840000.0ns 0V 303320000.0ns 0V 303360000.0ns 0.13183090090751648V 304080000.0ns 0.13183090090751648V 304120000.0ns 0.13183090090751648V 304600000.0ns 0.13183090090751648V 304640000.0ns 0.13183090090751648V 305360000.0ns 0.13183090090751648V 305400000.0ns 0.13183090090751648V 305880000.0ns 0.13183090090751648V 305920000.0ns 0.13183090090751648V 306640000.0ns 0.13183090090751648V 306680000.0ns 0V 307160000.0ns 0V 307200000.0ns 0.2884390950202942V 307920000.0ns 0.2884390950202942V 307960000.0ns 0.2884390950202942V 308440000.0ns 0.2884390950202942V 308480000.0ns 0.2884390950202942V 309200000.0ns 0.2884390950202942V 309240000.0ns 0.2884390950202942V 309720000.0ns 0.2884390950202942V 309760000.0ns 0.2884390950202942V 310480000.0ns 0.2884390950202942V 310520000.0ns 0V 311000000.0ns 0V 311040000.0ns 0.28828611969947815V 311760000.0ns 0.28828611969947815V 311800000.0ns 0.28828611969947815V 312280000.0ns 0.28828611969947815V 312320000.0ns 0.28828611969947815V 313040000.0ns 0.28828611969947815V 313080000.0ns 0.28828611969947815V 313560000.0ns 0.28828611969947815V 313600000.0ns 0.28828611969947815V 314320000.0ns 0.28828611969947815V 314360000.0ns 0V 314840000.0ns 0V 314880000.0ns 0.12186630815267563V 315600000.0ns 0.12186630815267563V 315640000.0ns 0.12186630815267563V 316120000.0ns 0.12186630815267563V 316160000.0ns 0.12186630815267563V 316880000.0ns 0.12186630815267563V 316920000.0ns 0.12186630815267563V 317400000.0ns 0.12186630815267563V 317440000.0ns 0.12186630815267563V 318160000.0ns 0.12186630815267563V 318200000.0ns 0V 318680000.0ns 0V 318720000.0ns 0.19145509600639343V 319440000.0ns 0.19145509600639343V 319480000.0ns 0.19145509600639343V 319960000.0ns 0.19145509600639343V 320000000.0ns 0.19145509600639343V 320720000.0ns 0.19145509600639343V 320760000.0ns 0.19145509600639343V 321240000.0ns 0.19145509600639343V 321280000.0ns 0.19145509600639343V 322000000.0ns 0.19145509600639343V 322040000.0ns 0V 322520000.0ns 0V 322560000.0ns 0.11054428666830063V 323280000.0ns 0.11054428666830063V 323320000.0ns 0.11054428666830063V 323800000.0ns 0.11054428666830063V 323840000.0ns 0.11054428666830063V 324560000.0ns 0.11054428666830063V 324600000.0ns 0.11054428666830063V 325080000.0ns 0.11054428666830063V 325120000.0ns 0.11054428666830063V 325840000.0ns 0.11054428666830063V 325880000.0ns 0V 326360000.0ns 0V 326400000.0ns 0.21930380165576935V 327120000.0ns 0.21930380165576935V 327160000.0ns 0.21930380165576935V 327640000.0ns 0.21930380165576935V 327680000.0ns 0.21930380165576935V 328400000.0ns 0.21930380165576935V 328440000.0ns 0.21930380165576935V 328920000.0ns 0.21930380165576935V 328960000.0ns 0.21930380165576935V 329680000.0ns 0.21930380165576935V 329720000.0ns 0V 330200000.0ns 0V 330240000.0ns 0.2989511489868164V 330960000.0ns 0.2989511489868164V 331000000.0ns 0.2989511489868164V 331480000.0ns 0.2989511489868164V 331520000.0ns 0.2989511489868164V 332240000.0ns 0.2989511489868164V 332280000.0ns 0.2989511489868164V 332760000.0ns 0.2989511489868164V 332800000.0ns 0.2989511489868164V 333520000.0ns 0.2989511489868164V 333560000.0ns 0V 334040000.0ns 0V 334080000.0ns 0.1375253051519394V 334800000.0ns 0.1375253051519394V 334840000.0ns 0.1375253051519394V 335320000.0ns 0.1375253051519394V 335360000.0ns 0.1375253051519394V 336080000.0ns 0.1375253051519394V 336120000.0ns 0.1375253051519394V 336600000.0ns 0.1375253051519394V 336640000.0ns 0.1375253051519394V 337360000.0ns 0.1375253051519394V 337400000.0ns 0V 337880000.0ns 0V 337920000.0ns 0.22864295542240143V 338640000.0ns 0.22864295542240143V 338680000.0ns 0.22864295542240143V 339160000.0ns 0.22864295542240143V 339200000.0ns 0.22864295542240143V 339920000.0ns 0.22864295542240143V 339960000.0ns 0.22864295542240143V 340440000.0ns 0.22864295542240143V 340480000.0ns 0.22864295542240143V 341200000.0ns 0.22864295542240143V 341240000.0ns 0V 341720000.0ns 0V 341760000.0ns 0.2767345905303955V 342480000.0ns 0.2767345905303955V 342520000.0ns 0.2767345905303955V 343000000.0ns 0.2767345905303955V 343040000.0ns 0.2767345905303955V 343760000.0ns 0.2767345905303955V 343800000.0ns 0.2767345905303955V 344280000.0ns 0.2767345905303955V 344320000.0ns 0.2767345905303955V 345040000.0ns 0.2767345905303955V 345080000.0ns 0V 345560000.0ns 0V 345600000.0ns 0.28965499997138977V 346320000.0ns 0.28965499997138977V 346360000.0ns 0.28965499997138977V 346840000.0ns 0.28965499997138977V 346880000.0ns 0.28965499997138977V 347600000.0ns 0.28965499997138977V 347640000.0ns 0.28965499997138977V 348120000.0ns 0.28965499997138977V 348160000.0ns 0.28965499997138977V 348880000.0ns 0.28965499997138977V 348920000.0ns 0V 349400000.0ns 0V 349440000.0ns 0.11806777864694595V 350160000.0ns 0.11806777864694595V 350200000.0ns 0.11806777864694595V 350680000.0ns 0.11806777864694595V 350720000.0ns 0.11806777864694595V 351440000.0ns 0.11806777864694595V 351480000.0ns 0.11806777864694595V 351960000.0ns 0.11806777864694595V 352000000.0ns 0.11806777864694595V 352720000.0ns 0.11806777864694595V 352760000.0ns 0V 353240000.0ns 0V 353280000.0ns 0.29533690214157104V 354000000.0ns 0.29533690214157104V 354040000.0ns 0.29533690214157104V 354520000.0ns 0.29533690214157104V 354560000.0ns 0.29533690214157104V 355280000.0ns 0.29533690214157104V 355320000.0ns 0.29533690214157104V 355800000.0ns 0.29533690214157104V 355840000.0ns 0.29533690214157104V 356560000.0ns 0.29533690214157104V 356600000.0ns 0V 357080000.0ns 0V 357120000.0ns 0.2566644549369812V 357840000.0ns 0.2566644549369812V 357880000.0ns 0.2566644549369812V 358360000.0ns 0.2566644549369812V 358400000.0ns 0.2566644549369812V 359120000.0ns 0.2566644549369812V 359160000.0ns 0.2566644549369812V 359640000.0ns 0.2566644549369812V 359680000.0ns 0.2566644549369812V 360400000.0ns 0.2566644549369812V 360440000.0ns 0V 360920000.0ns 0V 360960000.0ns 0.24335122108459473V 361680000.0ns 0.24335122108459473V 361720000.0ns 0.24335122108459473V 362200000.0ns 0.24335122108459473V 362240000.0ns 0.24335122108459473V 362960000.0ns 0.24335122108459473V 363000000.0ns 0.24335122108459473V 363480000.0ns 0.24335122108459473V 363520000.0ns 0.24335122108459473V 364240000.0ns 0.24335122108459473V 364280000.0ns 0V 364760000.0ns 0V 364800000.0ns 0.10000113397836685V 365520000.0ns 0.10000113397836685V 365560000.0ns 0.10000113397836685V 366040000.0ns 0.10000113397836685V 366080000.0ns 0.10000113397836685V 366800000.0ns 0.10000113397836685V 366840000.0ns 0.10000113397836685V 367320000.0ns 0.10000113397836685V 367360000.0ns 0.10000113397836685V 368080000.0ns 0.10000113397836685V 368120000.0ns 0V 368600000.0ns 0V 368640000.0ns 0.29782530665397644V 369360000.0ns 0.29782530665397644V 369400000.0ns 0.29782530665397644V 369880000.0ns 0.29782530665397644V 369920000.0ns 0.29782530665397644V 370640000.0ns 0.29782530665397644V 370680000.0ns 0.29782530665397644V 371160000.0ns 0.29782530665397644V 371200000.0ns 0.29782530665397644V 371920000.0ns 0.29782530665397644V 371960000.0ns 0V 372440000.0ns 0V 372480000.0ns 0.15254473686218262V 373200000.0ns 0.15254473686218262V 373240000.0ns 0.15254473686218262V 373720000.0ns 0.15254473686218262V 373760000.0ns 0.15254473686218262V 374480000.0ns 0.15254473686218262V 374520000.0ns 0.15254473686218262V 375000000.0ns 0.15254473686218262V 375040000.0ns 0.15254473686218262V 375760000.0ns 0.15254473686218262V 375800000.0ns 0V 376280000.0ns 0V 376320000.0ns 0.1607566773891449V 377040000.0ns 0.1607566773891449V 377080000.0ns 0.1607566773891449V 377560000.0ns 0.1607566773891449V 377600000.0ns 0.1607566773891449V 378320000.0ns 0.1607566773891449V 378360000.0ns 0.1607566773891449V 378840000.0ns 0.1607566773891449V 378880000.0ns 0.1607566773891449V 379600000.0ns 0.1607566773891449V 379640000.0ns 0V 380120000.0ns 0V 380160000.0ns 0.13453927636146545V 380880000.0ns 0.13453927636146545V 380920000.0ns 0.13453927636146545V 381400000.0ns 0.13453927636146545V 381440000.0ns 0.13453927636146545V 382160000.0ns 0.13453927636146545V 382200000.0ns 0.13453927636146545V 382680000.0ns 0.13453927636146545V 382720000.0ns 0.13453927636146545V 383440000.0ns 0.13453927636146545V 383480000.0ns 0V 383960000.0ns 0V 384000000.0ns 0.20831502974033356V 384720000.0ns 0.20831502974033356V 384760000.0ns 0.20831502974033356V 385240000.0ns 0.20831502974033356V 385280000.0ns 0.20831502974033356V 386000000.0ns 0.20831502974033356V 386040000.0ns 0.20831502974033356V 386520000.0ns 0.20831502974033356V 386560000.0ns 0.20831502974033356V 387280000.0ns 0.20831502974033356V 387320000.0ns 0V 387800000.0ns 0V 387840000.0ns 0.2966122627258301V 388560000.0ns 0.2966122627258301V 388600000.0ns 0.2966122627258301V 389080000.0ns 0.2966122627258301V 389120000.0ns 0.2966122627258301V 389840000.0ns 0.2966122627258301V 389880000.0ns 0.2966122627258301V 390360000.0ns 0.2966122627258301V 390400000.0ns 0.2966122627258301V 391120000.0ns 0.2966122627258301V 391160000.0ns 0V)
BLOSS LOSS 0 v={(V(target_0)-V(Y_0)+V(Y_1))*(V(target_0)-V(Y_0)+V(Y_1))}
BNUDGE Y_0_NUDGED Y_1_NUDGED i={-1.0000000000000002e-06 * (V(target_0)-V(Y_0_FREE)+V(Y_1_FREE)) * V(NUDGED_OUTER)}
VVWWL_I0 WWL_I0 0 PWL(0ns 0V 40000.0ns 0V 80000.0ns 1.95V 480000.0ns 1.95V 520000.0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0V 8400000.0ns 0V 8440000.0ns 0V 8920000.0ns 0V 8960000.0ns 0V 9680000.0ns 0V 9720000.0ns 0V 10520000.0ns 0V 10560000.0ns 0V 10640000.0ns 0V 10680000.0ns 0V 11480000.0ns 0V 11520000.0ns 0V 12240000.0ns 0V 12280000.0ns 0V 12760000.0ns 0V 12800000.0ns 0V 13520000.0ns 0V 13560000.0ns 0V 14360000.0ns 0V 14400000.0ns 0V 14480000.0ns 0V 14520000.0ns 0V 15320000.0ns 0V 15360000.0ns 0V 16080000.0ns 0V 16120000.0ns 0V 16600000.0ns 0V 16640000.0ns 0V 17360000.0ns 0V 17400000.0ns 0V 18200000.0ns 0V 18240000.0ns 0V 18320000.0ns 0V 18360000.0ns 0V 19160000.0ns 0V 19200000.0ns 0V 19920000.0ns 0V 19960000.0ns 0V 20440000.0ns 0V 20480000.0ns 0V 21200000.0ns 0V 21240000.0ns 0V 22040000.0ns 0V 22080000.0ns 0V 22160000.0ns 0V 22200000.0ns 0V 23000000.0ns 0V 23040000.0ns 0V 23760000.0ns 0V 23800000.0ns 0V 24280000.0ns 0V 24320000.0ns 0V 25040000.0ns 0V 25080000.0ns 0V 25880000.0ns 0V 25920000.0ns 0V 26000000.0ns 0V 26040000.0ns 0V 26840000.0ns 0V 26880000.0ns 0V 27600000.0ns 0V 27640000.0ns 0V 28120000.0ns 0V 28160000.0ns 0V 28880000.0ns 0V 28920000.0ns 0V 29720000.0ns 0V 29760000.0ns 0V 29840000.0ns 0V 29880000.0ns 0V 30680000.0ns 0V 30720000.0ns 0V 31440000.0ns 0V 31480000.0ns 0V 31960000.0ns 0V 32000000.0ns 0V 32720000.0ns 0V 32760000.0ns 0V 33560000.0ns 0V 33600000.0ns 0V 33680000.0ns 0V 33720000.0ns 0V 34520000.0ns 0V 34560000.0ns 0V 35280000.0ns 0V 35320000.0ns 0V 35800000.0ns 0V 35840000.0ns 0V 36560000.0ns 0V 36600000.0ns 0V 37400000.0ns 0V 37440000.0ns 0V 37520000.0ns 0V 37560000.0ns 0V 38360000.0ns 0V 38400000.0ns 0V 39120000.0ns 0V 39160000.0ns 0V 39640000.0ns 0V 39680000.0ns 0V 40400000.0ns 0V 40440000.0ns 0V 41240000.0ns 0V 41280000.0ns 0V 41360000.0ns 0V 41400000.0ns 0V 42200000.0ns 0V 42240000.0ns 0V 42960000.0ns 0V 43000000.0ns 0V 43480000.0ns 0V 43520000.0ns 0V 44240000.0ns 0V 44280000.0ns 0V 45080000.0ns 0V 45120000.0ns 0V 45200000.0ns 0V 45240000.0ns 0V 46040000.0ns 0V 46080000.0ns 0V 46800000.0ns 0V 46840000.0ns 0V 47320000.0ns 0V 47360000.0ns 0V 48080000.0ns 0V 48120000.0ns 0V 48920000.0ns 0V 48960000.0ns 0V 49040000.0ns 0V 49080000.0ns 0V 49880000.0ns 0V 49920000.0ns 0V 50640000.0ns 0V 50680000.0ns 0V 51160000.0ns 0V 51200000.0ns 0V 51920000.0ns 0V 51960000.0ns 0V 52760000.0ns 0V 52800000.0ns 0V 52880000.0ns 0V 52920000.0ns 0V 53720000.0ns 0V 53760000.0ns 0V 54480000.0ns 0V 54520000.0ns 0V 55000000.0ns 0V 55040000.0ns 0V 55760000.0ns 0V 55800000.0ns 0V 56600000.0ns 0V 56640000.0ns 0V 56720000.0ns 0V 56760000.0ns 0V 57560000.0ns 0V 57600000.0ns 0V 58320000.0ns 0V 58360000.0ns 0V 58840000.0ns 0V 58880000.0ns 0V 59600000.0ns 0V 59640000.0ns 0V 60440000.0ns 0V 60480000.0ns 0V 60560000.0ns 0V 60600000.0ns 0V 61400000.0ns 0V 61440000.0ns 0V 62160000.0ns 0V 62200000.0ns 0V 62680000.0ns 0V 62720000.0ns 0V 63440000.0ns 0V 63480000.0ns 0V 64280000.0ns 0V 64320000.0ns 0V 64400000.0ns 0V 64440000.0ns 0V 65240000.0ns 0V 65280000.0ns 0V 66000000.0ns 0V 66040000.0ns 0V 66520000.0ns 0V 66560000.0ns 0V 67280000.0ns 0V 67320000.0ns 0V 68120000.0ns 0V 68160000.0ns 0V 68240000.0ns 0V 68280000.0ns 0V 69080000.0ns 0V 69120000.0ns 0V 69840000.0ns 0V 69880000.0ns 0V 70360000.0ns 0V 70400000.0ns 0V 71120000.0ns 0V 71160000.0ns 0V 71960000.0ns 0V 72000000.0ns 0V 72080000.0ns 0V 72120000.0ns 0V 72920000.0ns 0V 72960000.0ns 0V 73680000.0ns 0V 73720000.0ns 0V 74200000.0ns 0V 74240000.0ns 0V 74960000.0ns 0V 75000000.0ns 0V 75800000.0ns 0V 75840000.0ns 0V 75920000.0ns 0V 75960000.0ns 0V 76760000.0ns 0V 76800000.0ns 0V 77520000.0ns 0V 77560000.0ns 0V 78040000.0ns 0V 78080000.0ns 0V 78800000.0ns 0V 78840000.0ns 0V 79640000.0ns 0V 79680000.0ns 0V 79760000.0ns 0V 79800000.0ns 0V 80600000.0ns 0V 80640000.0ns 0V 81360000.0ns 0V 81400000.0ns 0V 81880000.0ns 0V 81920000.0ns 0V 82640000.0ns 0V 82680000.0ns 0V 83480000.0ns 0V 83520000.0ns 0V 83600000.0ns 0V 83640000.0ns 0V 84440000.0ns 0V 84480000.0ns 0V 85200000.0ns 0V 85240000.0ns 0V 85720000.0ns 0V 85760000.0ns 0V 86480000.0ns 0V 86520000.0ns 0V 87320000.0ns 0V 87360000.0ns 0V 87440000.0ns 0V 87480000.0ns 0V 88280000.0ns 0V 88320000.0ns 0V 89040000.0ns 0V 89080000.0ns 0V 89560000.0ns 0V 89600000.0ns 0V 90320000.0ns 0V 90360000.0ns 0V 91160000.0ns 0V 91200000.0ns 0V 91280000.0ns 0V 91320000.0ns 0V 92120000.0ns 0V 92160000.0ns 0V 92880000.0ns 0V 92920000.0ns 0V 93400000.0ns 0V 93440000.0ns 0V 94160000.0ns 0V 94200000.0ns 0V 95000000.0ns 0V 95040000.0ns 0V 95120000.0ns 0V 95160000.0ns 0V 95960000.0ns 0V 96000000.0ns 0V 96720000.0ns 0V 96760000.0ns 0V 97240000.0ns 0V 97280000.0ns 0V 98000000.0ns 0V 98040000.0ns 0V 98840000.0ns 0V 98880000.0ns 0V 98960000.0ns 0V 99000000.0ns 0V 99800000.0ns 0V 99840000.0ns 0V 100560000.0ns 0V 100600000.0ns 0V 101080000.0ns 0V 101120000.0ns 0V 101840000.0ns 0V 101880000.0ns 0V 102680000.0ns 0V 102720000.0ns 0V 102800000.0ns 0V 102840000.0ns 0V 103640000.0ns 0V 103680000.0ns 0V 104400000.0ns 0V 104440000.0ns 0V 104920000.0ns 0V 104960000.0ns 0V 105680000.0ns 0V 105720000.0ns 0V 106520000.0ns 0V 106560000.0ns 0V 106640000.0ns 0V 106680000.0ns 0V 107480000.0ns 0V 107520000.0ns 0V 108240000.0ns 0V 108280000.0ns 0V 108760000.0ns 0V 108800000.0ns 0V 109520000.0ns 0V 109560000.0ns 0V 110360000.0ns 0V 110400000.0ns 0V 110480000.0ns 0V 110520000.0ns 0V 111320000.0ns 0V 111360000.0ns 0V 112080000.0ns 0V 112120000.0ns 0V 112600000.0ns 0V 112640000.0ns 0V 113360000.0ns 0V 113400000.0ns 0V 114200000.0ns 0V 114240000.0ns 0V 114320000.0ns 0V 114360000.0ns 0V 115160000.0ns 0V 115200000.0ns 0V 115920000.0ns 0V 115960000.0ns 0V 116440000.0ns 0V 116480000.0ns 0V 117200000.0ns 0V 117240000.0ns 0V 118040000.0ns 0V 118080000.0ns 0V 118160000.0ns 0V 118200000.0ns 0V 119000000.0ns 0V 119040000.0ns 0V 119760000.0ns 0V 119800000.0ns 0V 120280000.0ns 0V 120320000.0ns 0V 121040000.0ns 0V 121080000.0ns 0V 121880000.0ns 0V 121920000.0ns 0V 122000000.0ns 0V 122040000.0ns 0V 122840000.0ns 0V 122880000.0ns 0V 123600000.0ns 0V 123640000.0ns 0V 124120000.0ns 0V 124160000.0ns 0V 124880000.0ns 0V 124920000.0ns 0V 125720000.0ns 0V 125760000.0ns 0V 125840000.0ns 0V 125880000.0ns 0V 126680000.0ns 0V 126720000.0ns 0V 127440000.0ns 0V 127480000.0ns 0V 127960000.0ns 0V 128000000.0ns 0V 128720000.0ns 0V 128760000.0ns 0V 129560000.0ns 0V 129600000.0ns 0V 129680000.0ns 0V 129720000.0ns 0V 130520000.0ns 0V 130560000.0ns 0V 131280000.0ns 0V 131320000.0ns 0V 131800000.0ns 0V 131840000.0ns 0V 132560000.0ns 0V 132600000.0ns 0V 133400000.0ns 0V 133440000.0ns 0V 133520000.0ns 0V 133560000.0ns 0V 134360000.0ns 0V 134400000.0ns 0V 135120000.0ns 0V 135160000.0ns 0V 135640000.0ns 0V 135680000.0ns 0V 136400000.0ns 0V 136440000.0ns 0V 137240000.0ns 0V 137280000.0ns 0V 137360000.0ns 0V 137400000.0ns 0V 138200000.0ns 0V 138240000.0ns 0V 138960000.0ns 0V 139000000.0ns 0V 139480000.0ns 0V 139520000.0ns 0V 140240000.0ns 0V 140280000.0ns 0V 141080000.0ns 0V 141120000.0ns 0V 141200000.0ns 0V 141240000.0ns 0V 142040000.0ns 0V 142080000.0ns 0V 142800000.0ns 0V 142840000.0ns 0V 143320000.0ns 0V 143360000.0ns 0V 144080000.0ns 0V 144120000.0ns 0V 144920000.0ns 0V 144960000.0ns 0V 145040000.0ns 0V 145080000.0ns 0V 145880000.0ns 0V 145920000.0ns 0V 146640000.0ns 0V 146680000.0ns 0V 147160000.0ns 0V 147200000.0ns 0V 147920000.0ns 0V 147960000.0ns 0V 148760000.0ns 0V 148800000.0ns 0V 148880000.0ns 0V 148920000.0ns 0V 149720000.0ns 0V 149760000.0ns 0V 150480000.0ns 0V 150520000.0ns 0V 151000000.0ns 0V 151040000.0ns 0V 151760000.0ns 0V 151800000.0ns 0V 152600000.0ns 0V 152640000.0ns 0V 152720000.0ns 0V 152760000.0ns 0V 153560000.0ns 0V 153600000.0ns 0V 154320000.0ns 0V 154360000.0ns 0V 154840000.0ns 0V 154880000.0ns 0V 155600000.0ns 0V 155640000.0ns 0V 156440000.0ns 0V 156480000.0ns 0V 156560000.0ns 0V 156600000.0ns 0V 157400000.0ns 0V 157440000.0ns 0V 158160000.0ns 0V 158200000.0ns 0V 158680000.0ns 0V 158720000.0ns 0V 159440000.0ns 0V 159480000.0ns 0V 160280000.0ns 0V 160320000.0ns 0V 160400000.0ns 0V 160440000.0ns 0V 161240000.0ns 0V 161280000.0ns 0V 162000000.0ns 0V 162040000.0ns 0V 162520000.0ns 0V 162560000.0ns 0V 163280000.0ns 0V 163320000.0ns 0V 164120000.0ns 0V 164160000.0ns 0V 164240000.0ns 0V 164280000.0ns 0V 165080000.0ns 0V 165120000.0ns 0V 165840000.0ns 0V 165880000.0ns 0V 166360000.0ns 0V 166400000.0ns 0V 167120000.0ns 0V 167160000.0ns 0V 167960000.0ns 0V 168000000.0ns 0V 168080000.0ns 0V 168120000.0ns 0V 168920000.0ns 0V 168960000.0ns 0V 169680000.0ns 0V 169720000.0ns 0V 170200000.0ns 0V 170240000.0ns 0V 170960000.0ns 0V 171000000.0ns 0V 171800000.0ns 0V 171840000.0ns 0V 171920000.0ns 0V 171960000.0ns 0V 172760000.0ns 0V 172800000.0ns 0V 173520000.0ns 0V 173560000.0ns 0V 174040000.0ns 0V 174080000.0ns 0V 174800000.0ns 0V 174840000.0ns 0V 175640000.0ns 0V 175680000.0ns 0V 175760000.0ns 0V 175800000.0ns 0V 176600000.0ns 0V 176640000.0ns 0V 177360000.0ns 0V 177400000.0ns 0V 177880000.0ns 0V 177920000.0ns 0V 178640000.0ns 0V 178680000.0ns 0V 179480000.0ns 0V 179520000.0ns 0V 179600000.0ns 0V 179640000.0ns 0V 180440000.0ns 0V 180480000.0ns 0V 181200000.0ns 0V 181240000.0ns 0V 181720000.0ns 0V 181760000.0ns 0V 182480000.0ns 0V 182520000.0ns 0V 183320000.0ns 0V 183360000.0ns 0V 183440000.0ns 0V 183480000.0ns 0V 184280000.0ns 0V 184320000.0ns 0V 185040000.0ns 0V 185080000.0ns 0V 185560000.0ns 0V 185600000.0ns 0V 186320000.0ns 0V 186360000.0ns 0V 187160000.0ns 0V 187200000.0ns 0V 187280000.0ns 0V 187320000.0ns 0V 188120000.0ns 0V 188160000.0ns 0V 188880000.0ns 0V 188920000.0ns 0V 189400000.0ns 0V 189440000.0ns 0V 190160000.0ns 0V 190200000.0ns 0V 191000000.0ns 0V 191040000.0ns 0V 191120000.0ns 0V 191160000.0ns 0V 191960000.0ns 0V 192000000.0ns 0V 192720000.0ns 0V 192760000.0ns 0V 193240000.0ns 0V 193280000.0ns 0V 194000000.0ns 0V 194040000.0ns 0V 194840000.0ns 0V 194880000.0ns 0V 194960000.0ns 0V 195000000.0ns 0V 195800000.0ns 0V 195840000.0ns 0V 196560000.0ns 0V 196600000.0ns 0V 197080000.0ns 0V 197120000.0ns 0V 197840000.0ns 0V 197880000.0ns 0V 198680000.0ns 0V 198720000.0ns 0V 198800000.0ns 0V 198840000.0ns 0V 199640000.0ns 0V 199680000.0ns 0V 200400000.0ns 0V 200440000.0ns 0V 200920000.0ns 0V 200960000.0ns 0V 201680000.0ns 0V 201720000.0ns 0V 202520000.0ns 0V 202560000.0ns 0V 202640000.0ns 0V 202680000.0ns 0V 203480000.0ns 0V 203520000.0ns 0V 204240000.0ns 0V 204280000.0ns 0V 204760000.0ns 0V 204800000.0ns 0V 205520000.0ns 0V 205560000.0ns 0V 206360000.0ns 0V 206400000.0ns 0V 206480000.0ns 0V 206520000.0ns 0V 207320000.0ns 0V 207360000.0ns 0V 208080000.0ns 0V 208120000.0ns 0V 208600000.0ns 0V 208640000.0ns 0V 209360000.0ns 0V 209400000.0ns 0V 210200000.0ns 0V 210240000.0ns 0V 210320000.0ns 0V 210360000.0ns 0V 211160000.0ns 0V 211200000.0ns 0V 211920000.0ns 0V 211960000.0ns 0V 212440000.0ns 0V 212480000.0ns 0V 213200000.0ns 0V 213240000.0ns 0V 214040000.0ns 0V 214080000.0ns 0V 214160000.0ns 0V 214200000.0ns 0V 215000000.0ns 0V 215040000.0ns 0V 215760000.0ns 0V 215800000.0ns 0V 216280000.0ns 0V 216320000.0ns 0V 217040000.0ns 0V 217080000.0ns 0V 217880000.0ns 0V 217920000.0ns 0V 218000000.0ns 0V 218040000.0ns 0V 218840000.0ns 0V 218880000.0ns 0V 219600000.0ns 0V 219640000.0ns 0V 220120000.0ns 0V 220160000.0ns 0V 220880000.0ns 0V 220920000.0ns 0V 221720000.0ns 0V 221760000.0ns 0V 221840000.0ns 0V 221880000.0ns 0V 222680000.0ns 0V 222720000.0ns 0V 223440000.0ns 0V 223480000.0ns 0V 223960000.0ns 0V 224000000.0ns 0V 224720000.0ns 0V 224760000.0ns 0V 225560000.0ns 0V 225600000.0ns 0V 225680000.0ns 0V 225720000.0ns 0V 226520000.0ns 0V 226560000.0ns 0V 227280000.0ns 0V 227320000.0ns 0V 227800000.0ns 0V 227840000.0ns 0V 228560000.0ns 0V 228600000.0ns 0V 229400000.0ns 0V 229440000.0ns 0V 229520000.0ns 0V 229560000.0ns 0V 230360000.0ns 0V 230400000.0ns 0V 231120000.0ns 0V 231160000.0ns 0V 231640000.0ns 0V 231680000.0ns 0V 232400000.0ns 0V 232440000.0ns 0V 233240000.0ns 0V 233280000.0ns 0V 233360000.0ns 0V 233400000.0ns 0V 234200000.0ns 0V 234240000.0ns 0V 234960000.0ns 0V 235000000.0ns 0V 235480000.0ns 0V 235520000.0ns 0V 236240000.0ns 0V 236280000.0ns 0V 237080000.0ns 0V 237120000.0ns 0V 237200000.0ns 0V 237240000.0ns 0V 238040000.0ns 0V 238080000.0ns 0V 238800000.0ns 0V 238840000.0ns 0V 239320000.0ns 0V 239360000.0ns 0V 240080000.0ns 0V 240120000.0ns 0V 240920000.0ns 0V 240960000.0ns 0V 241040000.0ns 0V 241080000.0ns 0V 241880000.0ns 0V 241920000.0ns 0V 242640000.0ns 0V 242680000.0ns 0V 243160000.0ns 0V 243200000.0ns 0V 243920000.0ns 0V 243960000.0ns 0V 244760000.0ns 0V 244800000.0ns 0V 244880000.0ns 0V 244920000.0ns 0V 245720000.0ns 0V 245760000.0ns 0V 246480000.0ns 0V 246520000.0ns 0V 247000000.0ns 0V 247040000.0ns 0V 247760000.0ns 0V 247800000.0ns 0V 248600000.0ns 0V 248640000.0ns 0V 248720000.0ns 0V 248760000.0ns 0V 249560000.0ns 0V 249600000.0ns 0V 250320000.0ns 0V 250360000.0ns 0V 250840000.0ns 0V 250880000.0ns 0V 251600000.0ns 0V 251640000.0ns 0V 252440000.0ns 0V 252480000.0ns 0V 252560000.0ns 0V 252600000.0ns 0V 253400000.0ns 0V 253440000.0ns 0V 254160000.0ns 0V 254200000.0ns 0V 254680000.0ns 0V 254720000.0ns 0V 255440000.0ns 0V 255480000.0ns 0V 256280000.0ns 0V 256320000.0ns 0V 256400000.0ns 0V 256440000.0ns 0V 257240000.0ns 0V 257280000.0ns 0V 258000000.0ns 0V 258040000.0ns 0V 258520000.0ns 0V 258560000.0ns 0V 259280000.0ns 0V 259320000.0ns 0V 260120000.0ns 0V 260160000.0ns 0V 260240000.0ns 0V 260280000.0ns 0V 261080000.0ns 0V 261120000.0ns 0V 261840000.0ns 0V 261880000.0ns 0V 262360000.0ns 0V 262400000.0ns 0V 263120000.0ns 0V 263160000.0ns 0V 263960000.0ns 0V 264000000.0ns 0V 264080000.0ns 0V 264120000.0ns 0V 264920000.0ns 0V 264960000.0ns 0V 265680000.0ns 0V 265720000.0ns 0V 266200000.0ns 0V 266240000.0ns 0V 266960000.0ns 0V 267000000.0ns 0V 267800000.0ns 0V 267840000.0ns 0V 267920000.0ns 0V 267960000.0ns 0V 268760000.0ns 0V 268800000.0ns 0V 269520000.0ns 0V 269560000.0ns 0V 270040000.0ns 0V 270080000.0ns 0V 270800000.0ns 0V 270840000.0ns 0V 271640000.0ns 0V 271680000.0ns 0V 271760000.0ns 0V 271800000.0ns 0V 272600000.0ns 0V 272640000.0ns 0V 273360000.0ns 0V 273400000.0ns 0V 273880000.0ns 0V 273920000.0ns 0V 274640000.0ns 0V 274680000.0ns 0V 275480000.0ns 0V 275520000.0ns 0V 275600000.0ns 0V 275640000.0ns 0V 276440000.0ns 0V 276480000.0ns 0V 277200000.0ns 0V 277240000.0ns 0V 277720000.0ns 0V 277760000.0ns 0V 278480000.0ns 0V 278520000.0ns 0V 279320000.0ns 0V 279360000.0ns 0V 279440000.0ns 0V 279480000.0ns 0V 280280000.0ns 0V 280320000.0ns 0V 281040000.0ns 0V 281080000.0ns 0V 281560000.0ns 0V 281600000.0ns 0V 282320000.0ns 0V 282360000.0ns 0V 283160000.0ns 0V 283200000.0ns 0V 283280000.0ns 0V 283320000.0ns 0V 284120000.0ns 0V 284160000.0ns 0V 284880000.0ns 0V 284920000.0ns 0V 285400000.0ns 0V 285440000.0ns 0V 286160000.0ns 0V 286200000.0ns 0V 287000000.0ns 0V 287040000.0ns 0V 287120000.0ns 0V 287160000.0ns 0V 287960000.0ns 0V 288000000.0ns 0V 288720000.0ns 0V 288760000.0ns 0V 289240000.0ns 0V 289280000.0ns 0V 290000000.0ns 0V 290040000.0ns 0V 290840000.0ns 0V 290880000.0ns 0V 290960000.0ns 0V 291000000.0ns 0V 291800000.0ns 0V 291840000.0ns 0V 292560000.0ns 0V 292600000.0ns 0V 293080000.0ns 0V 293120000.0ns 0V 293840000.0ns 0V 293880000.0ns 0V 294680000.0ns 0V 294720000.0ns 0V 294800000.0ns 0V 294840000.0ns 0V 295640000.0ns 0V 295680000.0ns 0V 296400000.0ns 0V 296440000.0ns 0V 296920000.0ns 0V 296960000.0ns 0V 297680000.0ns 0V 297720000.0ns 0V 298520000.0ns 0V 298560000.0ns 0V 298640000.0ns 0V 298680000.0ns 0V 299480000.0ns 0V 299520000.0ns 0V 300240000.0ns 0V 300280000.0ns 0V 300760000.0ns 0V 300800000.0ns 0V 301520000.0ns 0V 301560000.0ns 0V 302360000.0ns 0V 302400000.0ns 0V 302480000.0ns 0V 302520000.0ns 0V 303320000.0ns 0V 303360000.0ns 0V 304080000.0ns 0V 304120000.0ns 0V 304600000.0ns 0V 304640000.0ns 0V 305360000.0ns 0V 305400000.0ns 0V 306200000.0ns 0V 306240000.0ns 0V 306320000.0ns 0V 306360000.0ns 0V 307160000.0ns 0V 307200000.0ns 0V 307920000.0ns 0V 307960000.0ns 0V 308440000.0ns 0V 308480000.0ns 0V 309200000.0ns 0V 309240000.0ns 0V 310040000.0ns 0V 310080000.0ns 0V 310160000.0ns 0V 310200000.0ns 0V 311000000.0ns 0V 311040000.0ns 0V 311760000.0ns 0V 311800000.0ns 0V 312280000.0ns 0V 312320000.0ns 0V 313040000.0ns 0V 313080000.0ns 0V 313880000.0ns 0V 313920000.0ns 0V 314000000.0ns 0V 314040000.0ns 0V 314840000.0ns 0V 314880000.0ns 0V 315600000.0ns 0V 315640000.0ns 0V 316120000.0ns 0V 316160000.0ns 0V 316880000.0ns 0V 316920000.0ns 0V 317720000.0ns 0V 317760000.0ns 0V 317840000.0ns 0V 317880000.0ns 0V 318680000.0ns 0V 318720000.0ns 0V 319440000.0ns 0V 319480000.0ns 0V 319960000.0ns 0V 320000000.0ns 0V 320720000.0ns 0V 320760000.0ns 0V 321560000.0ns 0V 321600000.0ns 0V 321680000.0ns 0V 321720000.0ns 0V 322520000.0ns 0V 322560000.0ns 0V 323280000.0ns 0V 323320000.0ns 0V 323800000.0ns 0V 323840000.0ns 0V 324560000.0ns 0V 324600000.0ns 0V 325400000.0ns 0V 325440000.0ns 0V 325520000.0ns 0V 325560000.0ns 0V 326360000.0ns 0V 326400000.0ns 0V 327120000.0ns 0V 327160000.0ns 0V 327640000.0ns 0V 327680000.0ns 0V 328400000.0ns 0V 328440000.0ns 0V 329240000.0ns 0V 329280000.0ns 0V 329360000.0ns 0V 329400000.0ns 0V 330200000.0ns 0V 330240000.0ns 0V 330960000.0ns 0V 331000000.0ns 0V 331480000.0ns 0V 331520000.0ns 0V 332240000.0ns 0V 332280000.0ns 0V 333080000.0ns 0V 333120000.0ns 0V 333200000.0ns 0V 333240000.0ns 0V 334040000.0ns 0V 334080000.0ns 0V 334800000.0ns 0V 334840000.0ns 0V 335320000.0ns 0V 335360000.0ns 0V 336080000.0ns 0V 336120000.0ns 0V 336920000.0ns 0V 336960000.0ns 0V 337040000.0ns 0V 337080000.0ns 0V 337880000.0ns 0V 337920000.0ns 0V 338640000.0ns 0V 338680000.0ns 0V 339160000.0ns 0V 339200000.0ns 0V 339920000.0ns 0V 339960000.0ns 0V 340760000.0ns 0V 340800000.0ns 0V 340880000.0ns 0V 340920000.0ns 0V 341720000.0ns 0V 341760000.0ns 0V 342480000.0ns 0V 342520000.0ns 0V 343000000.0ns 0V 343040000.0ns 0V 343760000.0ns 0V 343800000.0ns 0V 344600000.0ns 0V 344640000.0ns 0V 344720000.0ns 0V 344760000.0ns 0V 345560000.0ns 0V 345600000.0ns 0V 346320000.0ns 0V 346360000.0ns 0V 346840000.0ns 0V 346880000.0ns 0V 347600000.0ns 0V 347640000.0ns 0V 348440000.0ns 0V 348480000.0ns 0V 348560000.0ns 0V 348600000.0ns 0V 349400000.0ns 0V 349440000.0ns 0V 350160000.0ns 0V 350200000.0ns 0V 350680000.0ns 0V 350720000.0ns 0V 351440000.0ns 0V 351480000.0ns 0V 352280000.0ns 0V 352320000.0ns 0V 352400000.0ns 0V 352440000.0ns 0V 353240000.0ns 0V 353280000.0ns 0V 354000000.0ns 0V 354040000.0ns 0V 354520000.0ns 0V 354560000.0ns 0V 355280000.0ns 0V 355320000.0ns 0V 356120000.0ns 0V 356160000.0ns 0V 356240000.0ns 0V 356280000.0ns 0V 357080000.0ns 0V 357120000.0ns 0V 357840000.0ns 0V 357880000.0ns 0V 358360000.0ns 0V 358400000.0ns 0V 359120000.0ns 0V 359160000.0ns 0V 359960000.0ns 0V 360000000.0ns 0V 360080000.0ns 0V 360120000.0ns 0V 360920000.0ns 0V 360960000.0ns 0V 361680000.0ns 0V 361720000.0ns 0V 362200000.0ns 0V 362240000.0ns 0V 362960000.0ns 0V 363000000.0ns 0V 363800000.0ns 0V 363840000.0ns 0V 363920000.0ns 0V 363960000.0ns 0V 364760000.0ns 0V 364800000.0ns 0V 365520000.0ns 0V 365560000.0ns 0V 366040000.0ns 0V 366080000.0ns 0V 366800000.0ns 0V 366840000.0ns 0V 367640000.0ns 0V 367680000.0ns 0V 367760000.0ns 0V 367800000.0ns 0V 368600000.0ns 0V 368640000.0ns 0V 369360000.0ns 0V 369400000.0ns 0V 369880000.0ns 0V 369920000.0ns 0V 370640000.0ns 0V 370680000.0ns 0V 371480000.0ns 0V 371520000.0ns 0V 371600000.0ns 0V 371640000.0ns 0V 372440000.0ns 0V 372480000.0ns 0V 373200000.0ns 0V 373240000.0ns 0V 373720000.0ns 0V 373760000.0ns 0V 374480000.0ns 0V 374520000.0ns 0V 375320000.0ns 0V 375360000.0ns 0V 375440000.0ns 0V 375480000.0ns 0V 376280000.0ns 0V 376320000.0ns 0V 377040000.0ns 0V 377080000.0ns 0V 377560000.0ns 0V 377600000.0ns 0V 378320000.0ns 0V 378360000.0ns 0V 379160000.0ns 0V 379200000.0ns 0V 379280000.0ns 0V 379320000.0ns 0V 380120000.0ns 0V 380160000.0ns 0V 380880000.0ns 0V 380920000.0ns 0V 381400000.0ns 0V 381440000.0ns 0V 382160000.0ns 0V 382200000.0ns 0V 383000000.0ns 0V 383040000.0ns 0V 383120000.0ns 0V 383160000.0ns 0V 383960000.0ns 0V 384000000.0ns 0V 384720000.0ns 0V 384760000.0ns 0V 385240000.0ns 0V 385280000.0ns 0V 386000000.0ns 0V 386040000.0ns 0V 386840000.0ns 0V 386880000.0ns 0V 386960000.0ns 0V 387000000.0ns 0V 387800000.0ns 0V 387840000.0ns 0V 388560000.0ns 0V 388600000.0ns 0V 389080000.0ns 0V 389120000.0ns 0V 389840000.0ns 0V 389880000.0ns 0V 390680000.0ns 0V 390720000.0ns 0V 390800000.0ns 0V 390840000.0ns 0V)
VVWWL_J0 WWL_J0 0 PWL(0ns 0V 40000.0ns 0V 80000.0ns 1.95V 480000.0ns 1.95V 520000.0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0V 8400000.0ns 0V 8440000.0ns 0V 8920000.0ns 0V 8960000.0ns 0V 9680000.0ns 0V 9720000.0ns 0V 10520000.0ns 0V 10560000.0ns 0V 10640000.0ns 0V 10680000.0ns 0V 11480000.0ns 0V 11520000.0ns 0V 12240000.0ns 0V 12280000.0ns 0V 12760000.0ns 0V 12800000.0ns 0V 13520000.0ns 0V 13560000.0ns 0V 14360000.0ns 0V 14400000.0ns 0V 14480000.0ns 0V 14520000.0ns 0V 15320000.0ns 0V 15360000.0ns 0V 16080000.0ns 0V 16120000.0ns 0V 16600000.0ns 0V 16640000.0ns 0V 17360000.0ns 0V 17400000.0ns 0V 18200000.0ns 0V 18240000.0ns 0V 18320000.0ns 0V 18360000.0ns 0V 19160000.0ns 0V 19200000.0ns 0V 19920000.0ns 0V 19960000.0ns 0V 20440000.0ns 0V 20480000.0ns 0V 21200000.0ns 0V 21240000.0ns 0V 22040000.0ns 0V 22080000.0ns 0V 22160000.0ns 0V 22200000.0ns 0V 23000000.0ns 0V 23040000.0ns 0V 23760000.0ns 0V 23800000.0ns 0V 24280000.0ns 0V 24320000.0ns 0V 25040000.0ns 0V 25080000.0ns 0V 25880000.0ns 0V 25920000.0ns 0V 26000000.0ns 0V 26040000.0ns 0V 26840000.0ns 0V 26880000.0ns 0V 27600000.0ns 0V 27640000.0ns 0V 28120000.0ns 0V 28160000.0ns 0V 28880000.0ns 0V 28920000.0ns 0V 29720000.0ns 0V 29760000.0ns 0V 29840000.0ns 0V 29880000.0ns 0V 30680000.0ns 0V 30720000.0ns 0V 31440000.0ns 0V 31480000.0ns 0V 31960000.0ns 0V 32000000.0ns 0V 32720000.0ns 0V 32760000.0ns 0V 33560000.0ns 0V 33600000.0ns 0V 33680000.0ns 0V 33720000.0ns 0V 34520000.0ns 0V 34560000.0ns 0V 35280000.0ns 0V 35320000.0ns 0V 35800000.0ns 0V 35840000.0ns 0V 36560000.0ns 0V 36600000.0ns 0V 37400000.0ns 0V 37440000.0ns 0V 37520000.0ns 0V 37560000.0ns 0V 38360000.0ns 0V 38400000.0ns 0V 39120000.0ns 0V 39160000.0ns 0V 39640000.0ns 0V 39680000.0ns 0V 40400000.0ns 0V 40440000.0ns 0V 41240000.0ns 0V 41280000.0ns 0V 41360000.0ns 0V 41400000.0ns 0V 42200000.0ns 0V 42240000.0ns 0V 42960000.0ns 0V 43000000.0ns 0V 43480000.0ns 0V 43520000.0ns 0V 44240000.0ns 0V 44280000.0ns 0V 45080000.0ns 0V 45120000.0ns 0V 45200000.0ns 0V 45240000.0ns 0V 46040000.0ns 0V 46080000.0ns 0V 46800000.0ns 0V 46840000.0ns 0V 47320000.0ns 0V 47360000.0ns 0V 48080000.0ns 0V 48120000.0ns 0V 48920000.0ns 0V 48960000.0ns 0V 49040000.0ns 0V 49080000.0ns 0V 49880000.0ns 0V 49920000.0ns 0V 50640000.0ns 0V 50680000.0ns 0V 51160000.0ns 0V 51200000.0ns 0V 51920000.0ns 0V 51960000.0ns 0V 52760000.0ns 0V 52800000.0ns 0V 52880000.0ns 0V 52920000.0ns 0V 53720000.0ns 0V 53760000.0ns 0V 54480000.0ns 0V 54520000.0ns 0V 55000000.0ns 0V 55040000.0ns 0V 55760000.0ns 0V 55800000.0ns 0V 56600000.0ns 0V 56640000.0ns 0V 56720000.0ns 0V 56760000.0ns 0V 57560000.0ns 0V 57600000.0ns 0V 58320000.0ns 0V 58360000.0ns 0V 58840000.0ns 0V 58880000.0ns 0V 59600000.0ns 0V 59640000.0ns 0V 60440000.0ns 0V 60480000.0ns 0V 60560000.0ns 0V 60600000.0ns 0V 61400000.0ns 0V 61440000.0ns 0V 62160000.0ns 0V 62200000.0ns 0V 62680000.0ns 0V 62720000.0ns 0V 63440000.0ns 0V 63480000.0ns 0V 64280000.0ns 0V 64320000.0ns 0V 64400000.0ns 0V 64440000.0ns 0V 65240000.0ns 0V 65280000.0ns 0V 66000000.0ns 0V 66040000.0ns 0V 66520000.0ns 0V 66560000.0ns 0V 67280000.0ns 0V 67320000.0ns 0V 68120000.0ns 0V 68160000.0ns 0V 68240000.0ns 0V 68280000.0ns 0V 69080000.0ns 0V 69120000.0ns 0V 69840000.0ns 0V 69880000.0ns 0V 70360000.0ns 0V 70400000.0ns 0V 71120000.0ns 0V 71160000.0ns 0V 71960000.0ns 0V 72000000.0ns 0V 72080000.0ns 0V 72120000.0ns 0V 72920000.0ns 0V 72960000.0ns 0V 73680000.0ns 0V 73720000.0ns 0V 74200000.0ns 0V 74240000.0ns 0V 74960000.0ns 0V 75000000.0ns 0V 75800000.0ns 0V 75840000.0ns 0V 75920000.0ns 0V 75960000.0ns 0V 76760000.0ns 0V 76800000.0ns 0V 77520000.0ns 0V 77560000.0ns 0V 78040000.0ns 0V 78080000.0ns 0V 78800000.0ns 0V 78840000.0ns 0V 79640000.0ns 0V 79680000.0ns 0V 79760000.0ns 0V 79800000.0ns 0V 80600000.0ns 0V 80640000.0ns 0V 81360000.0ns 0V 81400000.0ns 0V 81880000.0ns 0V 81920000.0ns 0V 82640000.0ns 0V 82680000.0ns 0V 83480000.0ns 0V 83520000.0ns 0V 83600000.0ns 0V 83640000.0ns 0V 84440000.0ns 0V 84480000.0ns 0V 85200000.0ns 0V 85240000.0ns 0V 85720000.0ns 0V 85760000.0ns 0V 86480000.0ns 0V 86520000.0ns 0V 87320000.0ns 0V 87360000.0ns 0V 87440000.0ns 0V 87480000.0ns 0V 88280000.0ns 0V 88320000.0ns 0V 89040000.0ns 0V 89080000.0ns 0V 89560000.0ns 0V 89600000.0ns 0V 90320000.0ns 0V 90360000.0ns 0V 91160000.0ns 0V 91200000.0ns 0V 91280000.0ns 0V 91320000.0ns 0V 92120000.0ns 0V 92160000.0ns 0V 92880000.0ns 0V 92920000.0ns 0V 93400000.0ns 0V 93440000.0ns 0V 94160000.0ns 0V 94200000.0ns 0V 95000000.0ns 0V 95040000.0ns 0V 95120000.0ns 0V 95160000.0ns 0V 95960000.0ns 0V 96000000.0ns 0V 96720000.0ns 0V 96760000.0ns 0V 97240000.0ns 0V 97280000.0ns 0V 98000000.0ns 0V 98040000.0ns 0V 98840000.0ns 0V 98880000.0ns 0V 98960000.0ns 0V 99000000.0ns 0V 99800000.0ns 0V 99840000.0ns 0V 100560000.0ns 0V 100600000.0ns 0V 101080000.0ns 0V 101120000.0ns 0V 101840000.0ns 0V 101880000.0ns 0V 102680000.0ns 0V 102720000.0ns 0V 102800000.0ns 0V 102840000.0ns 0V 103640000.0ns 0V 103680000.0ns 0V 104400000.0ns 0V 104440000.0ns 0V 104920000.0ns 0V 104960000.0ns 0V 105680000.0ns 0V 105720000.0ns 0V 106520000.0ns 0V 106560000.0ns 0V 106640000.0ns 0V 106680000.0ns 0V 107480000.0ns 0V 107520000.0ns 0V 108240000.0ns 0V 108280000.0ns 0V 108760000.0ns 0V 108800000.0ns 0V 109520000.0ns 0V 109560000.0ns 0V 110360000.0ns 0V 110400000.0ns 0V 110480000.0ns 0V 110520000.0ns 0V 111320000.0ns 0V 111360000.0ns 0V 112080000.0ns 0V 112120000.0ns 0V 112600000.0ns 0V 112640000.0ns 0V 113360000.0ns 0V 113400000.0ns 0V 114200000.0ns 0V 114240000.0ns 0V 114320000.0ns 0V 114360000.0ns 0V 115160000.0ns 0V 115200000.0ns 0V 115920000.0ns 0V 115960000.0ns 0V 116440000.0ns 0V 116480000.0ns 0V 117200000.0ns 0V 117240000.0ns 0V 118040000.0ns 0V 118080000.0ns 0V 118160000.0ns 0V 118200000.0ns 0V 119000000.0ns 0V 119040000.0ns 0V 119760000.0ns 0V 119800000.0ns 0V 120280000.0ns 0V 120320000.0ns 0V 121040000.0ns 0V 121080000.0ns 0V 121880000.0ns 0V 121920000.0ns 0V 122000000.0ns 0V 122040000.0ns 0V 122840000.0ns 0V 122880000.0ns 0V 123600000.0ns 0V 123640000.0ns 0V 124120000.0ns 0V 124160000.0ns 0V 124880000.0ns 0V 124920000.0ns 0V 125720000.0ns 0V 125760000.0ns 0V 125840000.0ns 0V 125880000.0ns 0V 126680000.0ns 0V 126720000.0ns 0V 127440000.0ns 0V 127480000.0ns 0V 127960000.0ns 0V 128000000.0ns 0V 128720000.0ns 0V 128760000.0ns 0V 129560000.0ns 0V 129600000.0ns 0V 129680000.0ns 0V 129720000.0ns 0V 130520000.0ns 0V 130560000.0ns 0V 131280000.0ns 0V 131320000.0ns 0V 131800000.0ns 0V 131840000.0ns 0V 132560000.0ns 0V 132600000.0ns 0V 133400000.0ns 0V 133440000.0ns 0V 133520000.0ns 0V 133560000.0ns 0V 134360000.0ns 0V 134400000.0ns 0V 135120000.0ns 0V 135160000.0ns 0V 135640000.0ns 0V 135680000.0ns 0V 136400000.0ns 0V 136440000.0ns 0V 137240000.0ns 0V 137280000.0ns 0V 137360000.0ns 0V 137400000.0ns 0V 138200000.0ns 0V 138240000.0ns 0V 138960000.0ns 0V 139000000.0ns 0V 139480000.0ns 0V 139520000.0ns 0V 140240000.0ns 0V 140280000.0ns 0V 141080000.0ns 0V 141120000.0ns 0V 141200000.0ns 0V 141240000.0ns 0V 142040000.0ns 0V 142080000.0ns 0V 142800000.0ns 0V 142840000.0ns 0V 143320000.0ns 0V 143360000.0ns 0V 144080000.0ns 0V 144120000.0ns 0V 144920000.0ns 0V 144960000.0ns 0V 145040000.0ns 0V 145080000.0ns 0V 145880000.0ns 0V 145920000.0ns 0V 146640000.0ns 0V 146680000.0ns 0V 147160000.0ns 0V 147200000.0ns 0V 147920000.0ns 0V 147960000.0ns 0V 148760000.0ns 0V 148800000.0ns 0V 148880000.0ns 0V 148920000.0ns 0V 149720000.0ns 0V 149760000.0ns 0V 150480000.0ns 0V 150520000.0ns 0V 151000000.0ns 0V 151040000.0ns 0V 151760000.0ns 0V 151800000.0ns 0V 152600000.0ns 0V 152640000.0ns 0V 152720000.0ns 0V 152760000.0ns 0V 153560000.0ns 0V 153600000.0ns 0V 154320000.0ns 0V 154360000.0ns 0V 154840000.0ns 0V 154880000.0ns 0V 155600000.0ns 0V 155640000.0ns 0V 156440000.0ns 0V 156480000.0ns 0V 156560000.0ns 0V 156600000.0ns 0V 157400000.0ns 0V 157440000.0ns 0V 158160000.0ns 0V 158200000.0ns 0V 158680000.0ns 0V 158720000.0ns 0V 159440000.0ns 0V 159480000.0ns 0V 160280000.0ns 0V 160320000.0ns 0V 160400000.0ns 0V 160440000.0ns 0V 161240000.0ns 0V 161280000.0ns 0V 162000000.0ns 0V 162040000.0ns 0V 162520000.0ns 0V 162560000.0ns 0V 163280000.0ns 0V 163320000.0ns 0V 164120000.0ns 0V 164160000.0ns 0V 164240000.0ns 0V 164280000.0ns 0V 165080000.0ns 0V 165120000.0ns 0V 165840000.0ns 0V 165880000.0ns 0V 166360000.0ns 0V 166400000.0ns 0V 167120000.0ns 0V 167160000.0ns 0V 167960000.0ns 0V 168000000.0ns 0V 168080000.0ns 0V 168120000.0ns 0V 168920000.0ns 0V 168960000.0ns 0V 169680000.0ns 0V 169720000.0ns 0V 170200000.0ns 0V 170240000.0ns 0V 170960000.0ns 0V 171000000.0ns 0V 171800000.0ns 0V 171840000.0ns 0V 171920000.0ns 0V 171960000.0ns 0V 172760000.0ns 0V 172800000.0ns 0V 173520000.0ns 0V 173560000.0ns 0V 174040000.0ns 0V 174080000.0ns 0V 174800000.0ns 0V 174840000.0ns 0V 175640000.0ns 0V 175680000.0ns 0V 175760000.0ns 0V 175800000.0ns 0V 176600000.0ns 0V 176640000.0ns 0V 177360000.0ns 0V 177400000.0ns 0V 177880000.0ns 0V 177920000.0ns 0V 178640000.0ns 0V 178680000.0ns 0V 179480000.0ns 0V 179520000.0ns 0V 179600000.0ns 0V 179640000.0ns 0V 180440000.0ns 0V 180480000.0ns 0V 181200000.0ns 0V 181240000.0ns 0V 181720000.0ns 0V 181760000.0ns 0V 182480000.0ns 0V 182520000.0ns 0V 183320000.0ns 0V 183360000.0ns 0V 183440000.0ns 0V 183480000.0ns 0V 184280000.0ns 0V 184320000.0ns 0V 185040000.0ns 0V 185080000.0ns 0V 185560000.0ns 0V 185600000.0ns 0V 186320000.0ns 0V 186360000.0ns 0V 187160000.0ns 0V 187200000.0ns 0V 187280000.0ns 0V 187320000.0ns 0V 188120000.0ns 0V 188160000.0ns 0V 188880000.0ns 0V 188920000.0ns 0V 189400000.0ns 0V 189440000.0ns 0V 190160000.0ns 0V 190200000.0ns 0V 191000000.0ns 0V 191040000.0ns 0V 191120000.0ns 0V 191160000.0ns 0V 191960000.0ns 0V 192000000.0ns 0V 192720000.0ns 0V 192760000.0ns 0V 193240000.0ns 0V 193280000.0ns 0V 194000000.0ns 0V 194040000.0ns 0V 194840000.0ns 0V 194880000.0ns 0V 194960000.0ns 0V 195000000.0ns 0V 195800000.0ns 0V 195840000.0ns 0V 196560000.0ns 0V 196600000.0ns 0V 197080000.0ns 0V 197120000.0ns 0V 197840000.0ns 0V 197880000.0ns 0V 198680000.0ns 0V 198720000.0ns 0V 198800000.0ns 0V 198840000.0ns 0V 199640000.0ns 0V 199680000.0ns 0V 200400000.0ns 0V 200440000.0ns 0V 200920000.0ns 0V 200960000.0ns 0V 201680000.0ns 0V 201720000.0ns 0V 202520000.0ns 0V 202560000.0ns 0V 202640000.0ns 0V 202680000.0ns 0V 203480000.0ns 0V 203520000.0ns 0V 204240000.0ns 0V 204280000.0ns 0V 204760000.0ns 0V 204800000.0ns 0V 205520000.0ns 0V 205560000.0ns 0V 206360000.0ns 0V 206400000.0ns 0V 206480000.0ns 0V 206520000.0ns 0V 207320000.0ns 0V 207360000.0ns 0V 208080000.0ns 0V 208120000.0ns 0V 208600000.0ns 0V 208640000.0ns 0V 209360000.0ns 0V 209400000.0ns 0V 210200000.0ns 0V 210240000.0ns 0V 210320000.0ns 0V 210360000.0ns 0V 211160000.0ns 0V 211200000.0ns 0V 211920000.0ns 0V 211960000.0ns 0V 212440000.0ns 0V 212480000.0ns 0V 213200000.0ns 0V 213240000.0ns 0V 214040000.0ns 0V 214080000.0ns 0V 214160000.0ns 0V 214200000.0ns 0V 215000000.0ns 0V 215040000.0ns 0V 215760000.0ns 0V 215800000.0ns 0V 216280000.0ns 0V 216320000.0ns 0V 217040000.0ns 0V 217080000.0ns 0V 217880000.0ns 0V 217920000.0ns 0V 218000000.0ns 0V 218040000.0ns 0V 218840000.0ns 0V 218880000.0ns 0V 219600000.0ns 0V 219640000.0ns 0V 220120000.0ns 0V 220160000.0ns 0V 220880000.0ns 0V 220920000.0ns 0V 221720000.0ns 0V 221760000.0ns 0V 221840000.0ns 0V 221880000.0ns 0V 222680000.0ns 0V 222720000.0ns 0V 223440000.0ns 0V 223480000.0ns 0V 223960000.0ns 0V 224000000.0ns 0V 224720000.0ns 0V 224760000.0ns 0V 225560000.0ns 0V 225600000.0ns 0V 225680000.0ns 0V 225720000.0ns 0V 226520000.0ns 0V 226560000.0ns 0V 227280000.0ns 0V 227320000.0ns 0V 227800000.0ns 0V 227840000.0ns 0V 228560000.0ns 0V 228600000.0ns 0V 229400000.0ns 0V 229440000.0ns 0V 229520000.0ns 0V 229560000.0ns 0V 230360000.0ns 0V 230400000.0ns 0V 231120000.0ns 0V 231160000.0ns 0V 231640000.0ns 0V 231680000.0ns 0V 232400000.0ns 0V 232440000.0ns 0V 233240000.0ns 0V 233280000.0ns 0V 233360000.0ns 0V 233400000.0ns 0V 234200000.0ns 0V 234240000.0ns 0V 234960000.0ns 0V 235000000.0ns 0V 235480000.0ns 0V 235520000.0ns 0V 236240000.0ns 0V 236280000.0ns 0V 237080000.0ns 0V 237120000.0ns 0V 237200000.0ns 0V 237240000.0ns 0V 238040000.0ns 0V 238080000.0ns 0V 238800000.0ns 0V 238840000.0ns 0V 239320000.0ns 0V 239360000.0ns 0V 240080000.0ns 0V 240120000.0ns 0V 240920000.0ns 0V 240960000.0ns 0V 241040000.0ns 0V 241080000.0ns 0V 241880000.0ns 0V 241920000.0ns 0V 242640000.0ns 0V 242680000.0ns 0V 243160000.0ns 0V 243200000.0ns 0V 243920000.0ns 0V 243960000.0ns 0V 244760000.0ns 0V 244800000.0ns 0V 244880000.0ns 0V 244920000.0ns 0V 245720000.0ns 0V 245760000.0ns 0V 246480000.0ns 0V 246520000.0ns 0V 247000000.0ns 0V 247040000.0ns 0V 247760000.0ns 0V 247800000.0ns 0V 248600000.0ns 0V 248640000.0ns 0V 248720000.0ns 0V 248760000.0ns 0V 249560000.0ns 0V 249600000.0ns 0V 250320000.0ns 0V 250360000.0ns 0V 250840000.0ns 0V 250880000.0ns 0V 251600000.0ns 0V 251640000.0ns 0V 252440000.0ns 0V 252480000.0ns 0V 252560000.0ns 0V 252600000.0ns 0V 253400000.0ns 0V 253440000.0ns 0V 254160000.0ns 0V 254200000.0ns 0V 254680000.0ns 0V 254720000.0ns 0V 255440000.0ns 0V 255480000.0ns 0V 256280000.0ns 0V 256320000.0ns 0V 256400000.0ns 0V 256440000.0ns 0V 257240000.0ns 0V 257280000.0ns 0V 258000000.0ns 0V 258040000.0ns 0V 258520000.0ns 0V 258560000.0ns 0V 259280000.0ns 0V 259320000.0ns 0V 260120000.0ns 0V 260160000.0ns 0V 260240000.0ns 0V 260280000.0ns 0V 261080000.0ns 0V 261120000.0ns 0V 261840000.0ns 0V 261880000.0ns 0V 262360000.0ns 0V 262400000.0ns 0V 263120000.0ns 0V 263160000.0ns 0V 263960000.0ns 0V 264000000.0ns 0V 264080000.0ns 0V 264120000.0ns 0V 264920000.0ns 0V 264960000.0ns 0V 265680000.0ns 0V 265720000.0ns 0V 266200000.0ns 0V 266240000.0ns 0V 266960000.0ns 0V 267000000.0ns 0V 267800000.0ns 0V 267840000.0ns 0V 267920000.0ns 0V 267960000.0ns 0V 268760000.0ns 0V 268800000.0ns 0V 269520000.0ns 0V 269560000.0ns 0V 270040000.0ns 0V 270080000.0ns 0V 270800000.0ns 0V 270840000.0ns 0V 271640000.0ns 0V 271680000.0ns 0V 271760000.0ns 0V 271800000.0ns 0V 272600000.0ns 0V 272640000.0ns 0V 273360000.0ns 0V 273400000.0ns 0V 273880000.0ns 0V 273920000.0ns 0V 274640000.0ns 0V 274680000.0ns 0V 275480000.0ns 0V 275520000.0ns 0V 275600000.0ns 0V 275640000.0ns 0V 276440000.0ns 0V 276480000.0ns 0V 277200000.0ns 0V 277240000.0ns 0V 277720000.0ns 0V 277760000.0ns 0V 278480000.0ns 0V 278520000.0ns 0V 279320000.0ns 0V 279360000.0ns 0V 279440000.0ns 0V 279480000.0ns 0V 280280000.0ns 0V 280320000.0ns 0V 281040000.0ns 0V 281080000.0ns 0V 281560000.0ns 0V 281600000.0ns 0V 282320000.0ns 0V 282360000.0ns 0V 283160000.0ns 0V 283200000.0ns 0V 283280000.0ns 0V 283320000.0ns 0V 284120000.0ns 0V 284160000.0ns 0V 284880000.0ns 0V 284920000.0ns 0V 285400000.0ns 0V 285440000.0ns 0V 286160000.0ns 0V 286200000.0ns 0V 287000000.0ns 0V 287040000.0ns 0V 287120000.0ns 0V 287160000.0ns 0V 287960000.0ns 0V 288000000.0ns 0V 288720000.0ns 0V 288760000.0ns 0V 289240000.0ns 0V 289280000.0ns 0V 290000000.0ns 0V 290040000.0ns 0V 290840000.0ns 0V 290880000.0ns 0V 290960000.0ns 0V 291000000.0ns 0V 291800000.0ns 0V 291840000.0ns 0V 292560000.0ns 0V 292600000.0ns 0V 293080000.0ns 0V 293120000.0ns 0V 293840000.0ns 0V 293880000.0ns 0V 294680000.0ns 0V 294720000.0ns 0V 294800000.0ns 0V 294840000.0ns 0V 295640000.0ns 0V 295680000.0ns 0V 296400000.0ns 0V 296440000.0ns 0V 296920000.0ns 0V 296960000.0ns 0V 297680000.0ns 0V 297720000.0ns 0V 298520000.0ns 0V 298560000.0ns 0V 298640000.0ns 0V 298680000.0ns 0V 299480000.0ns 0V 299520000.0ns 0V 300240000.0ns 0V 300280000.0ns 0V 300760000.0ns 0V 300800000.0ns 0V 301520000.0ns 0V 301560000.0ns 0V 302360000.0ns 0V 302400000.0ns 0V 302480000.0ns 0V 302520000.0ns 0V 303320000.0ns 0V 303360000.0ns 0V 304080000.0ns 0V 304120000.0ns 0V 304600000.0ns 0V 304640000.0ns 0V 305360000.0ns 0V 305400000.0ns 0V 306200000.0ns 0V 306240000.0ns 0V 306320000.0ns 0V 306360000.0ns 0V 307160000.0ns 0V 307200000.0ns 0V 307920000.0ns 0V 307960000.0ns 0V 308440000.0ns 0V 308480000.0ns 0V 309200000.0ns 0V 309240000.0ns 0V 310040000.0ns 0V 310080000.0ns 0V 310160000.0ns 0V 310200000.0ns 0V 311000000.0ns 0V 311040000.0ns 0V 311760000.0ns 0V 311800000.0ns 0V 312280000.0ns 0V 312320000.0ns 0V 313040000.0ns 0V 313080000.0ns 0V 313880000.0ns 0V 313920000.0ns 0V 314000000.0ns 0V 314040000.0ns 0V 314840000.0ns 0V 314880000.0ns 0V 315600000.0ns 0V 315640000.0ns 0V 316120000.0ns 0V 316160000.0ns 0V 316880000.0ns 0V 316920000.0ns 0V 317720000.0ns 0V 317760000.0ns 0V 317840000.0ns 0V 317880000.0ns 0V 318680000.0ns 0V 318720000.0ns 0V 319440000.0ns 0V 319480000.0ns 0V 319960000.0ns 0V 320000000.0ns 0V 320720000.0ns 0V 320760000.0ns 0V 321560000.0ns 0V 321600000.0ns 0V 321680000.0ns 0V 321720000.0ns 0V 322520000.0ns 0V 322560000.0ns 0V 323280000.0ns 0V 323320000.0ns 0V 323800000.0ns 0V 323840000.0ns 0V 324560000.0ns 0V 324600000.0ns 0V 325400000.0ns 0V 325440000.0ns 0V 325520000.0ns 0V 325560000.0ns 0V 326360000.0ns 0V 326400000.0ns 0V 327120000.0ns 0V 327160000.0ns 0V 327640000.0ns 0V 327680000.0ns 0V 328400000.0ns 0V 328440000.0ns 0V 329240000.0ns 0V 329280000.0ns 0V 329360000.0ns 0V 329400000.0ns 0V 330200000.0ns 0V 330240000.0ns 0V 330960000.0ns 0V 331000000.0ns 0V 331480000.0ns 0V 331520000.0ns 0V 332240000.0ns 0V 332280000.0ns 0V 333080000.0ns 0V 333120000.0ns 0V 333200000.0ns 0V 333240000.0ns 0V 334040000.0ns 0V 334080000.0ns 0V 334800000.0ns 0V 334840000.0ns 0V 335320000.0ns 0V 335360000.0ns 0V 336080000.0ns 0V 336120000.0ns 0V 336920000.0ns 0V 336960000.0ns 0V 337040000.0ns 0V 337080000.0ns 0V 337880000.0ns 0V 337920000.0ns 0V 338640000.0ns 0V 338680000.0ns 0V 339160000.0ns 0V 339200000.0ns 0V 339920000.0ns 0V 339960000.0ns 0V 340760000.0ns 0V 340800000.0ns 0V 340880000.0ns 0V 340920000.0ns 0V 341720000.0ns 0V 341760000.0ns 0V 342480000.0ns 0V 342520000.0ns 0V 343000000.0ns 0V 343040000.0ns 0V 343760000.0ns 0V 343800000.0ns 0V 344600000.0ns 0V 344640000.0ns 0V 344720000.0ns 0V 344760000.0ns 0V 345560000.0ns 0V 345600000.0ns 0V 346320000.0ns 0V 346360000.0ns 0V 346840000.0ns 0V 346880000.0ns 0V 347600000.0ns 0V 347640000.0ns 0V 348440000.0ns 0V 348480000.0ns 0V 348560000.0ns 0V 348600000.0ns 0V 349400000.0ns 0V 349440000.0ns 0V 350160000.0ns 0V 350200000.0ns 0V 350680000.0ns 0V 350720000.0ns 0V 351440000.0ns 0V 351480000.0ns 0V 352280000.0ns 0V 352320000.0ns 0V 352400000.0ns 0V 352440000.0ns 0V 353240000.0ns 0V 353280000.0ns 0V 354000000.0ns 0V 354040000.0ns 0V 354520000.0ns 0V 354560000.0ns 0V 355280000.0ns 0V 355320000.0ns 0V 356120000.0ns 0V 356160000.0ns 0V 356240000.0ns 0V 356280000.0ns 0V 357080000.0ns 0V 357120000.0ns 0V 357840000.0ns 0V 357880000.0ns 0V 358360000.0ns 0V 358400000.0ns 0V 359120000.0ns 0V 359160000.0ns 0V 359960000.0ns 0V 360000000.0ns 0V 360080000.0ns 0V 360120000.0ns 0V 360920000.0ns 0V 360960000.0ns 0V 361680000.0ns 0V 361720000.0ns 0V 362200000.0ns 0V 362240000.0ns 0V 362960000.0ns 0V 363000000.0ns 0V 363800000.0ns 0V 363840000.0ns 0V 363920000.0ns 0V 363960000.0ns 0V 364760000.0ns 0V 364800000.0ns 0V 365520000.0ns 0V 365560000.0ns 0V 366040000.0ns 0V 366080000.0ns 0V 366800000.0ns 0V 366840000.0ns 0V 367640000.0ns 0V 367680000.0ns 0V 367760000.0ns 0V 367800000.0ns 0V 368600000.0ns 0V 368640000.0ns 0V 369360000.0ns 0V 369400000.0ns 0V 369880000.0ns 0V 369920000.0ns 0V 370640000.0ns 0V 370680000.0ns 0V 371480000.0ns 0V 371520000.0ns 0V 371600000.0ns 0V 371640000.0ns 0V 372440000.0ns 0V 372480000.0ns 0V 373200000.0ns 0V 373240000.0ns 0V 373720000.0ns 0V 373760000.0ns 0V 374480000.0ns 0V 374520000.0ns 0V 375320000.0ns 0V 375360000.0ns 0V 375440000.0ns 0V 375480000.0ns 0V 376280000.0ns 0V 376320000.0ns 0V 377040000.0ns 0V 377080000.0ns 0V 377560000.0ns 0V 377600000.0ns 0V 378320000.0ns 0V 378360000.0ns 0V 379160000.0ns 0V 379200000.0ns 0V 379280000.0ns 0V 379320000.0ns 0V 380120000.0ns 0V 380160000.0ns 0V 380880000.0ns 0V 380920000.0ns 0V 381400000.0ns 0V 381440000.0ns 0V 382160000.0ns 0V 382200000.0ns 0V 383000000.0ns 0V 383040000.0ns 0V 383120000.0ns 0V 383160000.0ns 0V 383960000.0ns 0V 384000000.0ns 0V 384720000.0ns 0V 384760000.0ns 0V 385240000.0ns 0V 385280000.0ns 0V 386000000.0ns 0V 386040000.0ns 0V 386840000.0ns 0V 386880000.0ns 0V 386960000.0ns 0V 387000000.0ns 0V 387800000.0ns 0V 387840000.0ns 0V 388560000.0ns 0V 388600000.0ns 0V 389080000.0ns 0V 389120000.0ns 0V 389840000.0ns 0V 389880000.0ns 0V 390680000.0ns 0V 390720000.0ns 0V 390800000.0ns 0V 390840000.0ns 0V)
VVWWL_I1 WWL_I1 0 PWL(0ns 0V 920000.0ns 0V 960000.0ns 1.95V 1360000.0ns 1.95V 1400000.0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0V 8400000.0ns 0V 8440000.0ns 0V 8920000.0ns 0V 8960000.0ns 0V 9680000.0ns 0V 9720000.0ns 0V 10520000.0ns 0V 10560000.0ns 0V 10640000.0ns 0V 10680000.0ns 0V 11480000.0ns 0V 11520000.0ns 0V 12240000.0ns 0V 12280000.0ns 0V 12760000.0ns 0V 12800000.0ns 0V 13520000.0ns 0V 13560000.0ns 0V 14360000.0ns 0V 14400000.0ns 0V 14480000.0ns 0V 14520000.0ns 0V 15320000.0ns 0V 15360000.0ns 0V 16080000.0ns 0V 16120000.0ns 0V 16600000.0ns 0V 16640000.0ns 0V 17360000.0ns 0V 17400000.0ns 0V 18200000.0ns 0V 18240000.0ns 0V 18320000.0ns 0V 18360000.0ns 0V 19160000.0ns 0V 19200000.0ns 0V 19920000.0ns 0V 19960000.0ns 0V 20440000.0ns 0V 20480000.0ns 0V 21200000.0ns 0V 21240000.0ns 0V 22040000.0ns 0V 22080000.0ns 0V 22160000.0ns 0V 22200000.0ns 0V 23000000.0ns 0V 23040000.0ns 0V 23760000.0ns 0V 23800000.0ns 0V 24280000.0ns 0V 24320000.0ns 0V 25040000.0ns 0V 25080000.0ns 0V 25880000.0ns 0V 25920000.0ns 0V 26000000.0ns 0V 26040000.0ns 0V 26840000.0ns 0V 26880000.0ns 0V 27600000.0ns 0V 27640000.0ns 0V 28120000.0ns 0V 28160000.0ns 0V 28880000.0ns 0V 28920000.0ns 0V 29720000.0ns 0V 29760000.0ns 0V 29840000.0ns 0V 29880000.0ns 0V 30680000.0ns 0V 30720000.0ns 0V 31440000.0ns 0V 31480000.0ns 0V 31960000.0ns 0V 32000000.0ns 0V 32720000.0ns 0V 32760000.0ns 0V 33560000.0ns 0V 33600000.0ns 0V 33680000.0ns 0V 33720000.0ns 0V 34520000.0ns 0V 34560000.0ns 0V 35280000.0ns 0V 35320000.0ns 0V 35800000.0ns 0V 35840000.0ns 0V 36560000.0ns 0V 36600000.0ns 0V 37400000.0ns 0V 37440000.0ns 0V 37520000.0ns 0V 37560000.0ns 0V 38360000.0ns 0V 38400000.0ns 0V 39120000.0ns 0V 39160000.0ns 0V 39640000.0ns 0V 39680000.0ns 0V 40400000.0ns 0V 40440000.0ns 0V 41240000.0ns 0V 41280000.0ns 0V 41360000.0ns 0V 41400000.0ns 0V 42200000.0ns 0V 42240000.0ns 0V 42960000.0ns 0V 43000000.0ns 0V 43480000.0ns 0V 43520000.0ns 0V 44240000.0ns 0V 44280000.0ns 0V 45080000.0ns 0V 45120000.0ns 0V 45200000.0ns 0V 45240000.0ns 0V 46040000.0ns 0V 46080000.0ns 0V 46800000.0ns 0V 46840000.0ns 0V 47320000.0ns 0V 47360000.0ns 0V 48080000.0ns 0V 48120000.0ns 0V 48920000.0ns 0V 48960000.0ns 0V 49040000.0ns 0V 49080000.0ns 0V 49880000.0ns 0V 49920000.0ns 0V 50640000.0ns 0V 50680000.0ns 0V 51160000.0ns 0V 51200000.0ns 0V 51920000.0ns 0V 51960000.0ns 0V 52760000.0ns 0V 52800000.0ns 0V 52880000.0ns 0V 52920000.0ns 0V 53720000.0ns 0V 53760000.0ns 0V 54480000.0ns 0V 54520000.0ns 0V 55000000.0ns 0V 55040000.0ns 0V 55760000.0ns 0V 55800000.0ns 0V 56600000.0ns 0V 56640000.0ns 0V 56720000.0ns 0V 56760000.0ns 0V 57560000.0ns 0V 57600000.0ns 0V 58320000.0ns 0V 58360000.0ns 0V 58840000.0ns 0V 58880000.0ns 0V 59600000.0ns 0V 59640000.0ns 0V 60440000.0ns 0V 60480000.0ns 0V 60560000.0ns 0V 60600000.0ns 0V 61400000.0ns 0V 61440000.0ns 0V 62160000.0ns 0V 62200000.0ns 0V 62680000.0ns 0V 62720000.0ns 0V 63440000.0ns 0V 63480000.0ns 0V 64280000.0ns 0V 64320000.0ns 0V 64400000.0ns 0V 64440000.0ns 0V 65240000.0ns 0V 65280000.0ns 0V 66000000.0ns 0V 66040000.0ns 0V 66520000.0ns 0V 66560000.0ns 0V 67280000.0ns 0V 67320000.0ns 0V 68120000.0ns 0V 68160000.0ns 0V 68240000.0ns 0V 68280000.0ns 0V 69080000.0ns 0V 69120000.0ns 0V 69840000.0ns 0V 69880000.0ns 0V 70360000.0ns 0V 70400000.0ns 0V 71120000.0ns 0V 71160000.0ns 0V 71960000.0ns 0V 72000000.0ns 0V 72080000.0ns 0V 72120000.0ns 0V 72920000.0ns 0V 72960000.0ns 0V 73680000.0ns 0V 73720000.0ns 0V 74200000.0ns 0V 74240000.0ns 0V 74960000.0ns 0V 75000000.0ns 0V 75800000.0ns 0V 75840000.0ns 0V 75920000.0ns 0V 75960000.0ns 0V 76760000.0ns 0V 76800000.0ns 0V 77520000.0ns 0V 77560000.0ns 0V 78040000.0ns 0V 78080000.0ns 0V 78800000.0ns 0V 78840000.0ns 0V 79640000.0ns 0V 79680000.0ns 0V 79760000.0ns 0V 79800000.0ns 0V 80600000.0ns 0V 80640000.0ns 0V 81360000.0ns 0V 81400000.0ns 0V 81880000.0ns 0V 81920000.0ns 0V 82640000.0ns 0V 82680000.0ns 0V 83480000.0ns 0V 83520000.0ns 0V 83600000.0ns 0V 83640000.0ns 0V 84440000.0ns 0V 84480000.0ns 0V 85200000.0ns 0V 85240000.0ns 0V 85720000.0ns 0V 85760000.0ns 0V 86480000.0ns 0V 86520000.0ns 0V 87320000.0ns 0V 87360000.0ns 0V 87440000.0ns 0V 87480000.0ns 0V 88280000.0ns 0V 88320000.0ns 0V 89040000.0ns 0V 89080000.0ns 0V 89560000.0ns 0V 89600000.0ns 0V 90320000.0ns 0V 90360000.0ns 0V 91160000.0ns 0V 91200000.0ns 0V 91280000.0ns 0V 91320000.0ns 0V 92120000.0ns 0V 92160000.0ns 0V 92880000.0ns 0V 92920000.0ns 0V 93400000.0ns 0V 93440000.0ns 0V 94160000.0ns 0V 94200000.0ns 0V 95000000.0ns 0V 95040000.0ns 0V 95120000.0ns 0V 95160000.0ns 0V 95960000.0ns 0V 96000000.0ns 0V 96720000.0ns 0V 96760000.0ns 0V 97240000.0ns 0V 97280000.0ns 0V 98000000.0ns 0V 98040000.0ns 0V 98840000.0ns 0V 98880000.0ns 0V 98960000.0ns 0V 99000000.0ns 0V 99800000.0ns 0V 99840000.0ns 0V 100560000.0ns 0V 100600000.0ns 0V 101080000.0ns 0V 101120000.0ns 0V 101840000.0ns 0V 101880000.0ns 0V 102680000.0ns 0V 102720000.0ns 0V 102800000.0ns 0V 102840000.0ns 0V 103640000.0ns 0V 103680000.0ns 0V 104400000.0ns 0V 104440000.0ns 0V 104920000.0ns 0V 104960000.0ns 0V 105680000.0ns 0V 105720000.0ns 0V 106520000.0ns 0V 106560000.0ns 0V 106640000.0ns 0V 106680000.0ns 0V 107480000.0ns 0V 107520000.0ns 0V 108240000.0ns 0V 108280000.0ns 0V 108760000.0ns 0V 108800000.0ns 0V 109520000.0ns 0V 109560000.0ns 0V 110360000.0ns 0V 110400000.0ns 0V 110480000.0ns 0V 110520000.0ns 0V 111320000.0ns 0V 111360000.0ns 0V 112080000.0ns 0V 112120000.0ns 0V 112600000.0ns 0V 112640000.0ns 0V 113360000.0ns 0V 113400000.0ns 0V 114200000.0ns 0V 114240000.0ns 0V 114320000.0ns 0V 114360000.0ns 0V 115160000.0ns 0V 115200000.0ns 0V 115920000.0ns 0V 115960000.0ns 0V 116440000.0ns 0V 116480000.0ns 0V 117200000.0ns 0V 117240000.0ns 0V 118040000.0ns 0V 118080000.0ns 0V 118160000.0ns 0V 118200000.0ns 0V 119000000.0ns 0V 119040000.0ns 0V 119760000.0ns 0V 119800000.0ns 0V 120280000.0ns 0V 120320000.0ns 0V 121040000.0ns 0V 121080000.0ns 0V 121880000.0ns 0V 121920000.0ns 0V 122000000.0ns 0V 122040000.0ns 0V 122840000.0ns 0V 122880000.0ns 0V 123600000.0ns 0V 123640000.0ns 0V 124120000.0ns 0V 124160000.0ns 0V 124880000.0ns 0V 124920000.0ns 0V 125720000.0ns 0V 125760000.0ns 0V 125840000.0ns 0V 125880000.0ns 0V 126680000.0ns 0V 126720000.0ns 0V 127440000.0ns 0V 127480000.0ns 0V 127960000.0ns 0V 128000000.0ns 0V 128720000.0ns 0V 128760000.0ns 0V 129560000.0ns 0V 129600000.0ns 0V 129680000.0ns 0V 129720000.0ns 0V 130520000.0ns 0V 130560000.0ns 0V 131280000.0ns 0V 131320000.0ns 0V 131800000.0ns 0V 131840000.0ns 0V 132560000.0ns 0V 132600000.0ns 0V 133400000.0ns 0V 133440000.0ns 0V 133520000.0ns 0V 133560000.0ns 0V 134360000.0ns 0V 134400000.0ns 0V 135120000.0ns 0V 135160000.0ns 0V 135640000.0ns 0V 135680000.0ns 0V 136400000.0ns 0V 136440000.0ns 0V 137240000.0ns 0V 137280000.0ns 0V 137360000.0ns 0V 137400000.0ns 0V 138200000.0ns 0V 138240000.0ns 0V 138960000.0ns 0V 139000000.0ns 0V 139480000.0ns 0V 139520000.0ns 0V 140240000.0ns 0V 140280000.0ns 0V 141080000.0ns 0V 141120000.0ns 0V 141200000.0ns 0V 141240000.0ns 0V 142040000.0ns 0V 142080000.0ns 0V 142800000.0ns 0V 142840000.0ns 0V 143320000.0ns 0V 143360000.0ns 0V 144080000.0ns 0V 144120000.0ns 0V 144920000.0ns 0V 144960000.0ns 0V 145040000.0ns 0V 145080000.0ns 0V 145880000.0ns 0V 145920000.0ns 0V 146640000.0ns 0V 146680000.0ns 0V 147160000.0ns 0V 147200000.0ns 0V 147920000.0ns 0V 147960000.0ns 0V 148760000.0ns 0V 148800000.0ns 0V 148880000.0ns 0V 148920000.0ns 0V 149720000.0ns 0V 149760000.0ns 0V 150480000.0ns 0V 150520000.0ns 0V 151000000.0ns 0V 151040000.0ns 0V 151760000.0ns 0V 151800000.0ns 0V 152600000.0ns 0V 152640000.0ns 0V 152720000.0ns 0V 152760000.0ns 0V 153560000.0ns 0V 153600000.0ns 0V 154320000.0ns 0V 154360000.0ns 0V 154840000.0ns 0V 154880000.0ns 0V 155600000.0ns 0V 155640000.0ns 0V 156440000.0ns 0V 156480000.0ns 0V 156560000.0ns 0V 156600000.0ns 0V 157400000.0ns 0V 157440000.0ns 0V 158160000.0ns 0V 158200000.0ns 0V 158680000.0ns 0V 158720000.0ns 0V 159440000.0ns 0V 159480000.0ns 0V 160280000.0ns 0V 160320000.0ns 0V 160400000.0ns 0V 160440000.0ns 0V 161240000.0ns 0V 161280000.0ns 0V 162000000.0ns 0V 162040000.0ns 0V 162520000.0ns 0V 162560000.0ns 0V 163280000.0ns 0V 163320000.0ns 0V 164120000.0ns 0V 164160000.0ns 0V 164240000.0ns 0V 164280000.0ns 0V 165080000.0ns 0V 165120000.0ns 0V 165840000.0ns 0V 165880000.0ns 0V 166360000.0ns 0V 166400000.0ns 0V 167120000.0ns 0V 167160000.0ns 0V 167960000.0ns 0V 168000000.0ns 0V 168080000.0ns 0V 168120000.0ns 0V 168920000.0ns 0V 168960000.0ns 0V 169680000.0ns 0V 169720000.0ns 0V 170200000.0ns 0V 170240000.0ns 0V 170960000.0ns 0V 171000000.0ns 0V 171800000.0ns 0V 171840000.0ns 0V 171920000.0ns 0V 171960000.0ns 0V 172760000.0ns 0V 172800000.0ns 0V 173520000.0ns 0V 173560000.0ns 0V 174040000.0ns 0V 174080000.0ns 0V 174800000.0ns 0V 174840000.0ns 0V 175640000.0ns 0V 175680000.0ns 0V 175760000.0ns 0V 175800000.0ns 0V 176600000.0ns 0V 176640000.0ns 0V 177360000.0ns 0V 177400000.0ns 0V 177880000.0ns 0V 177920000.0ns 0V 178640000.0ns 0V 178680000.0ns 0V 179480000.0ns 0V 179520000.0ns 0V 179600000.0ns 0V 179640000.0ns 0V 180440000.0ns 0V 180480000.0ns 0V 181200000.0ns 0V 181240000.0ns 0V 181720000.0ns 0V 181760000.0ns 0V 182480000.0ns 0V 182520000.0ns 0V 183320000.0ns 0V 183360000.0ns 0V 183440000.0ns 0V 183480000.0ns 0V 184280000.0ns 0V 184320000.0ns 0V 185040000.0ns 0V 185080000.0ns 0V 185560000.0ns 0V 185600000.0ns 0V 186320000.0ns 0V 186360000.0ns 0V 187160000.0ns 0V 187200000.0ns 0V 187280000.0ns 0V 187320000.0ns 0V 188120000.0ns 0V 188160000.0ns 0V 188880000.0ns 0V 188920000.0ns 0V 189400000.0ns 0V 189440000.0ns 0V 190160000.0ns 0V 190200000.0ns 0V 191000000.0ns 0V 191040000.0ns 0V 191120000.0ns 0V 191160000.0ns 0V 191960000.0ns 0V 192000000.0ns 0V 192720000.0ns 0V 192760000.0ns 0V 193240000.0ns 0V 193280000.0ns 0V 194000000.0ns 0V 194040000.0ns 0V 194840000.0ns 0V 194880000.0ns 0V 194960000.0ns 0V 195000000.0ns 0V 195800000.0ns 0V 195840000.0ns 0V 196560000.0ns 0V 196600000.0ns 0V 197080000.0ns 0V 197120000.0ns 0V 197840000.0ns 0V 197880000.0ns 0V 198680000.0ns 0V 198720000.0ns 0V 198800000.0ns 0V 198840000.0ns 0V 199640000.0ns 0V 199680000.0ns 0V 200400000.0ns 0V 200440000.0ns 0V 200920000.0ns 0V 200960000.0ns 0V 201680000.0ns 0V 201720000.0ns 0V 202520000.0ns 0V 202560000.0ns 0V 202640000.0ns 0V 202680000.0ns 0V 203480000.0ns 0V 203520000.0ns 0V 204240000.0ns 0V 204280000.0ns 0V 204760000.0ns 0V 204800000.0ns 0V 205520000.0ns 0V 205560000.0ns 0V 206360000.0ns 0V 206400000.0ns 0V 206480000.0ns 0V 206520000.0ns 0V 207320000.0ns 0V 207360000.0ns 0V 208080000.0ns 0V 208120000.0ns 0V 208600000.0ns 0V 208640000.0ns 0V 209360000.0ns 0V 209400000.0ns 0V 210200000.0ns 0V 210240000.0ns 0V 210320000.0ns 0V 210360000.0ns 0V 211160000.0ns 0V 211200000.0ns 0V 211920000.0ns 0V 211960000.0ns 0V 212440000.0ns 0V 212480000.0ns 0V 213200000.0ns 0V 213240000.0ns 0V 214040000.0ns 0V 214080000.0ns 0V 214160000.0ns 0V 214200000.0ns 0V 215000000.0ns 0V 215040000.0ns 0V 215760000.0ns 0V 215800000.0ns 0V 216280000.0ns 0V 216320000.0ns 0V 217040000.0ns 0V 217080000.0ns 0V 217880000.0ns 0V 217920000.0ns 0V 218000000.0ns 0V 218040000.0ns 0V 218840000.0ns 0V 218880000.0ns 0V 219600000.0ns 0V 219640000.0ns 0V 220120000.0ns 0V 220160000.0ns 0V 220880000.0ns 0V 220920000.0ns 0V 221720000.0ns 0V 221760000.0ns 0V 221840000.0ns 0V 221880000.0ns 0V 222680000.0ns 0V 222720000.0ns 0V 223440000.0ns 0V 223480000.0ns 0V 223960000.0ns 0V 224000000.0ns 0V 224720000.0ns 0V 224760000.0ns 0V 225560000.0ns 0V 225600000.0ns 0V 225680000.0ns 0V 225720000.0ns 0V 226520000.0ns 0V 226560000.0ns 0V 227280000.0ns 0V 227320000.0ns 0V 227800000.0ns 0V 227840000.0ns 0V 228560000.0ns 0V 228600000.0ns 0V 229400000.0ns 0V 229440000.0ns 0V 229520000.0ns 0V 229560000.0ns 0V 230360000.0ns 0V 230400000.0ns 0V 231120000.0ns 0V 231160000.0ns 0V 231640000.0ns 0V 231680000.0ns 0V 232400000.0ns 0V 232440000.0ns 0V 233240000.0ns 0V 233280000.0ns 0V 233360000.0ns 0V 233400000.0ns 0V 234200000.0ns 0V 234240000.0ns 0V 234960000.0ns 0V 235000000.0ns 0V 235480000.0ns 0V 235520000.0ns 0V 236240000.0ns 0V 236280000.0ns 0V 237080000.0ns 0V 237120000.0ns 0V 237200000.0ns 0V 237240000.0ns 0V 238040000.0ns 0V 238080000.0ns 0V 238800000.0ns 0V 238840000.0ns 0V 239320000.0ns 0V 239360000.0ns 0V 240080000.0ns 0V 240120000.0ns 0V 240920000.0ns 0V 240960000.0ns 0V 241040000.0ns 0V 241080000.0ns 0V 241880000.0ns 0V 241920000.0ns 0V 242640000.0ns 0V 242680000.0ns 0V 243160000.0ns 0V 243200000.0ns 0V 243920000.0ns 0V 243960000.0ns 0V 244760000.0ns 0V 244800000.0ns 0V 244880000.0ns 0V 244920000.0ns 0V 245720000.0ns 0V 245760000.0ns 0V 246480000.0ns 0V 246520000.0ns 0V 247000000.0ns 0V 247040000.0ns 0V 247760000.0ns 0V 247800000.0ns 0V 248600000.0ns 0V 248640000.0ns 0V 248720000.0ns 0V 248760000.0ns 0V 249560000.0ns 0V 249600000.0ns 0V 250320000.0ns 0V 250360000.0ns 0V 250840000.0ns 0V 250880000.0ns 0V 251600000.0ns 0V 251640000.0ns 0V 252440000.0ns 0V 252480000.0ns 0V 252560000.0ns 0V 252600000.0ns 0V 253400000.0ns 0V 253440000.0ns 0V 254160000.0ns 0V 254200000.0ns 0V 254680000.0ns 0V 254720000.0ns 0V 255440000.0ns 0V 255480000.0ns 0V 256280000.0ns 0V 256320000.0ns 0V 256400000.0ns 0V 256440000.0ns 0V 257240000.0ns 0V 257280000.0ns 0V 258000000.0ns 0V 258040000.0ns 0V 258520000.0ns 0V 258560000.0ns 0V 259280000.0ns 0V 259320000.0ns 0V 260120000.0ns 0V 260160000.0ns 0V 260240000.0ns 0V 260280000.0ns 0V 261080000.0ns 0V 261120000.0ns 0V 261840000.0ns 0V 261880000.0ns 0V 262360000.0ns 0V 262400000.0ns 0V 263120000.0ns 0V 263160000.0ns 0V 263960000.0ns 0V 264000000.0ns 0V 264080000.0ns 0V 264120000.0ns 0V 264920000.0ns 0V 264960000.0ns 0V 265680000.0ns 0V 265720000.0ns 0V 266200000.0ns 0V 266240000.0ns 0V 266960000.0ns 0V 267000000.0ns 0V 267800000.0ns 0V 267840000.0ns 0V 267920000.0ns 0V 267960000.0ns 0V 268760000.0ns 0V 268800000.0ns 0V 269520000.0ns 0V 269560000.0ns 0V 270040000.0ns 0V 270080000.0ns 0V 270800000.0ns 0V 270840000.0ns 0V 271640000.0ns 0V 271680000.0ns 0V 271760000.0ns 0V 271800000.0ns 0V 272600000.0ns 0V 272640000.0ns 0V 273360000.0ns 0V 273400000.0ns 0V 273880000.0ns 0V 273920000.0ns 0V 274640000.0ns 0V 274680000.0ns 0V 275480000.0ns 0V 275520000.0ns 0V 275600000.0ns 0V 275640000.0ns 0V 276440000.0ns 0V 276480000.0ns 0V 277200000.0ns 0V 277240000.0ns 0V 277720000.0ns 0V 277760000.0ns 0V 278480000.0ns 0V 278520000.0ns 0V 279320000.0ns 0V 279360000.0ns 0V 279440000.0ns 0V 279480000.0ns 0V 280280000.0ns 0V 280320000.0ns 0V 281040000.0ns 0V 281080000.0ns 0V 281560000.0ns 0V 281600000.0ns 0V 282320000.0ns 0V 282360000.0ns 0V 283160000.0ns 0V 283200000.0ns 0V 283280000.0ns 0V 283320000.0ns 0V 284120000.0ns 0V 284160000.0ns 0V 284880000.0ns 0V 284920000.0ns 0V 285400000.0ns 0V 285440000.0ns 0V 286160000.0ns 0V 286200000.0ns 0V 287000000.0ns 0V 287040000.0ns 0V 287120000.0ns 0V 287160000.0ns 0V 287960000.0ns 0V 288000000.0ns 0V 288720000.0ns 0V 288760000.0ns 0V 289240000.0ns 0V 289280000.0ns 0V 290000000.0ns 0V 290040000.0ns 0V 290840000.0ns 0V 290880000.0ns 0V 290960000.0ns 0V 291000000.0ns 0V 291800000.0ns 0V 291840000.0ns 0V 292560000.0ns 0V 292600000.0ns 0V 293080000.0ns 0V 293120000.0ns 0V 293840000.0ns 0V 293880000.0ns 0V 294680000.0ns 0V 294720000.0ns 0V 294800000.0ns 0V 294840000.0ns 0V 295640000.0ns 0V 295680000.0ns 0V 296400000.0ns 0V 296440000.0ns 0V 296920000.0ns 0V 296960000.0ns 0V 297680000.0ns 0V 297720000.0ns 0V 298520000.0ns 0V 298560000.0ns 0V 298640000.0ns 0V 298680000.0ns 0V 299480000.0ns 0V 299520000.0ns 0V 300240000.0ns 0V 300280000.0ns 0V 300760000.0ns 0V 300800000.0ns 0V 301520000.0ns 0V 301560000.0ns 0V 302360000.0ns 0V 302400000.0ns 0V 302480000.0ns 0V 302520000.0ns 0V 303320000.0ns 0V 303360000.0ns 0V 304080000.0ns 0V 304120000.0ns 0V 304600000.0ns 0V 304640000.0ns 0V 305360000.0ns 0V 305400000.0ns 0V 306200000.0ns 0V 306240000.0ns 0V 306320000.0ns 0V 306360000.0ns 0V 307160000.0ns 0V 307200000.0ns 0V 307920000.0ns 0V 307960000.0ns 0V 308440000.0ns 0V 308480000.0ns 0V 309200000.0ns 0V 309240000.0ns 0V 310040000.0ns 0V 310080000.0ns 0V 310160000.0ns 0V 310200000.0ns 0V 311000000.0ns 0V 311040000.0ns 0V 311760000.0ns 0V 311800000.0ns 0V 312280000.0ns 0V 312320000.0ns 0V 313040000.0ns 0V 313080000.0ns 0V 313880000.0ns 0V 313920000.0ns 0V 314000000.0ns 0V 314040000.0ns 0V 314840000.0ns 0V 314880000.0ns 0V 315600000.0ns 0V 315640000.0ns 0V 316120000.0ns 0V 316160000.0ns 0V 316880000.0ns 0V 316920000.0ns 0V 317720000.0ns 0V 317760000.0ns 0V 317840000.0ns 0V 317880000.0ns 0V 318680000.0ns 0V 318720000.0ns 0V 319440000.0ns 0V 319480000.0ns 0V 319960000.0ns 0V 320000000.0ns 0V 320720000.0ns 0V 320760000.0ns 0V 321560000.0ns 0V 321600000.0ns 0V 321680000.0ns 0V 321720000.0ns 0V 322520000.0ns 0V 322560000.0ns 0V 323280000.0ns 0V 323320000.0ns 0V 323800000.0ns 0V 323840000.0ns 0V 324560000.0ns 0V 324600000.0ns 0V 325400000.0ns 0V 325440000.0ns 0V 325520000.0ns 0V 325560000.0ns 0V 326360000.0ns 0V 326400000.0ns 0V 327120000.0ns 0V 327160000.0ns 0V 327640000.0ns 0V 327680000.0ns 0V 328400000.0ns 0V 328440000.0ns 0V 329240000.0ns 0V 329280000.0ns 0V 329360000.0ns 0V 329400000.0ns 0V 330200000.0ns 0V 330240000.0ns 0V 330960000.0ns 0V 331000000.0ns 0V 331480000.0ns 0V 331520000.0ns 0V 332240000.0ns 0V 332280000.0ns 0V 333080000.0ns 0V 333120000.0ns 0V 333200000.0ns 0V 333240000.0ns 0V 334040000.0ns 0V 334080000.0ns 0V 334800000.0ns 0V 334840000.0ns 0V 335320000.0ns 0V 335360000.0ns 0V 336080000.0ns 0V 336120000.0ns 0V 336920000.0ns 0V 336960000.0ns 0V 337040000.0ns 0V 337080000.0ns 0V 337880000.0ns 0V 337920000.0ns 0V 338640000.0ns 0V 338680000.0ns 0V 339160000.0ns 0V 339200000.0ns 0V 339920000.0ns 0V 339960000.0ns 0V 340760000.0ns 0V 340800000.0ns 0V 340880000.0ns 0V 340920000.0ns 0V 341720000.0ns 0V 341760000.0ns 0V 342480000.0ns 0V 342520000.0ns 0V 343000000.0ns 0V 343040000.0ns 0V 343760000.0ns 0V 343800000.0ns 0V 344600000.0ns 0V 344640000.0ns 0V 344720000.0ns 0V 344760000.0ns 0V 345560000.0ns 0V 345600000.0ns 0V 346320000.0ns 0V 346360000.0ns 0V 346840000.0ns 0V 346880000.0ns 0V 347600000.0ns 0V 347640000.0ns 0V 348440000.0ns 0V 348480000.0ns 0V 348560000.0ns 0V 348600000.0ns 0V 349400000.0ns 0V 349440000.0ns 0V 350160000.0ns 0V 350200000.0ns 0V 350680000.0ns 0V 350720000.0ns 0V 351440000.0ns 0V 351480000.0ns 0V 352280000.0ns 0V 352320000.0ns 0V 352400000.0ns 0V 352440000.0ns 0V 353240000.0ns 0V 353280000.0ns 0V 354000000.0ns 0V 354040000.0ns 0V 354520000.0ns 0V 354560000.0ns 0V 355280000.0ns 0V 355320000.0ns 0V 356120000.0ns 0V 356160000.0ns 0V 356240000.0ns 0V 356280000.0ns 0V 357080000.0ns 0V 357120000.0ns 0V 357840000.0ns 0V 357880000.0ns 0V 358360000.0ns 0V 358400000.0ns 0V 359120000.0ns 0V 359160000.0ns 0V 359960000.0ns 0V 360000000.0ns 0V 360080000.0ns 0V 360120000.0ns 0V 360920000.0ns 0V 360960000.0ns 0V 361680000.0ns 0V 361720000.0ns 0V 362200000.0ns 0V 362240000.0ns 0V 362960000.0ns 0V 363000000.0ns 0V 363800000.0ns 0V 363840000.0ns 0V 363920000.0ns 0V 363960000.0ns 0V 364760000.0ns 0V 364800000.0ns 0V 365520000.0ns 0V 365560000.0ns 0V 366040000.0ns 0V 366080000.0ns 0V 366800000.0ns 0V 366840000.0ns 0V 367640000.0ns 0V 367680000.0ns 0V 367760000.0ns 0V 367800000.0ns 0V 368600000.0ns 0V 368640000.0ns 0V 369360000.0ns 0V 369400000.0ns 0V 369880000.0ns 0V 369920000.0ns 0V 370640000.0ns 0V 370680000.0ns 0V 371480000.0ns 0V 371520000.0ns 0V 371600000.0ns 0V 371640000.0ns 0V 372440000.0ns 0V 372480000.0ns 0V 373200000.0ns 0V 373240000.0ns 0V 373720000.0ns 0V 373760000.0ns 0V 374480000.0ns 0V 374520000.0ns 0V 375320000.0ns 0V 375360000.0ns 0V 375440000.0ns 0V 375480000.0ns 0V 376280000.0ns 0V 376320000.0ns 0V 377040000.0ns 0V 377080000.0ns 0V 377560000.0ns 0V 377600000.0ns 0V 378320000.0ns 0V 378360000.0ns 0V 379160000.0ns 0V 379200000.0ns 0V 379280000.0ns 0V 379320000.0ns 0V 380120000.0ns 0V 380160000.0ns 0V 380880000.0ns 0V 380920000.0ns 0V 381400000.0ns 0V 381440000.0ns 0V 382160000.0ns 0V 382200000.0ns 0V 383000000.0ns 0V 383040000.0ns 0V 383120000.0ns 0V 383160000.0ns 0V 383960000.0ns 0V 384000000.0ns 0V 384720000.0ns 0V 384760000.0ns 0V 385240000.0ns 0V 385280000.0ns 0V 386000000.0ns 0V 386040000.0ns 0V 386840000.0ns 0V 386880000.0ns 0V 386960000.0ns 0V 387000000.0ns 0V 387800000.0ns 0V 387840000.0ns 0V 388560000.0ns 0V 388600000.0ns 0V 389080000.0ns 0V 389120000.0ns 0V 389840000.0ns 0V 389880000.0ns 0V 390680000.0ns 0V 390720000.0ns 0V 390800000.0ns 0V 390840000.0ns 0V)
VVWWL_J1 WWL_J1 0 PWL(0ns 0V 920000.0ns 0V 960000.0ns 1.95V 1360000.0ns 1.95V 1400000.0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0V 8400000.0ns 0V 8440000.0ns 0V 8920000.0ns 0V 8960000.0ns 0V 9680000.0ns 0V 9720000.0ns 0V 10520000.0ns 0V 10560000.0ns 0V 10640000.0ns 0V 10680000.0ns 0V 11480000.0ns 0V 11520000.0ns 0V 12240000.0ns 0V 12280000.0ns 0V 12760000.0ns 0V 12800000.0ns 0V 13520000.0ns 0V 13560000.0ns 0V 14360000.0ns 0V 14400000.0ns 0V 14480000.0ns 0V 14520000.0ns 0V 15320000.0ns 0V 15360000.0ns 0V 16080000.0ns 0V 16120000.0ns 0V 16600000.0ns 0V 16640000.0ns 0V 17360000.0ns 0V 17400000.0ns 0V 18200000.0ns 0V 18240000.0ns 0V 18320000.0ns 0V 18360000.0ns 0V 19160000.0ns 0V 19200000.0ns 0V 19920000.0ns 0V 19960000.0ns 0V 20440000.0ns 0V 20480000.0ns 0V 21200000.0ns 0V 21240000.0ns 0V 22040000.0ns 0V 22080000.0ns 0V 22160000.0ns 0V 22200000.0ns 0V 23000000.0ns 0V 23040000.0ns 0V 23760000.0ns 0V 23800000.0ns 0V 24280000.0ns 0V 24320000.0ns 0V 25040000.0ns 0V 25080000.0ns 0V 25880000.0ns 0V 25920000.0ns 0V 26000000.0ns 0V 26040000.0ns 0V 26840000.0ns 0V 26880000.0ns 0V 27600000.0ns 0V 27640000.0ns 0V 28120000.0ns 0V 28160000.0ns 0V 28880000.0ns 0V 28920000.0ns 0V 29720000.0ns 0V 29760000.0ns 0V 29840000.0ns 0V 29880000.0ns 0V 30680000.0ns 0V 30720000.0ns 0V 31440000.0ns 0V 31480000.0ns 0V 31960000.0ns 0V 32000000.0ns 0V 32720000.0ns 0V 32760000.0ns 0V 33560000.0ns 0V 33600000.0ns 0V 33680000.0ns 0V 33720000.0ns 0V 34520000.0ns 0V 34560000.0ns 0V 35280000.0ns 0V 35320000.0ns 0V 35800000.0ns 0V 35840000.0ns 0V 36560000.0ns 0V 36600000.0ns 0V 37400000.0ns 0V 37440000.0ns 0V 37520000.0ns 0V 37560000.0ns 0V 38360000.0ns 0V 38400000.0ns 0V 39120000.0ns 0V 39160000.0ns 0V 39640000.0ns 0V 39680000.0ns 0V 40400000.0ns 0V 40440000.0ns 0V 41240000.0ns 0V 41280000.0ns 0V 41360000.0ns 0V 41400000.0ns 0V 42200000.0ns 0V 42240000.0ns 0V 42960000.0ns 0V 43000000.0ns 0V 43480000.0ns 0V 43520000.0ns 0V 44240000.0ns 0V 44280000.0ns 0V 45080000.0ns 0V 45120000.0ns 0V 45200000.0ns 0V 45240000.0ns 0V 46040000.0ns 0V 46080000.0ns 0V 46800000.0ns 0V 46840000.0ns 0V 47320000.0ns 0V 47360000.0ns 0V 48080000.0ns 0V 48120000.0ns 0V 48920000.0ns 0V 48960000.0ns 0V 49040000.0ns 0V 49080000.0ns 0V 49880000.0ns 0V 49920000.0ns 0V 50640000.0ns 0V 50680000.0ns 0V 51160000.0ns 0V 51200000.0ns 0V 51920000.0ns 0V 51960000.0ns 0V 52760000.0ns 0V 52800000.0ns 0V 52880000.0ns 0V 52920000.0ns 0V 53720000.0ns 0V 53760000.0ns 0V 54480000.0ns 0V 54520000.0ns 0V 55000000.0ns 0V 55040000.0ns 0V 55760000.0ns 0V 55800000.0ns 0V 56600000.0ns 0V 56640000.0ns 0V 56720000.0ns 0V 56760000.0ns 0V 57560000.0ns 0V 57600000.0ns 0V 58320000.0ns 0V 58360000.0ns 0V 58840000.0ns 0V 58880000.0ns 0V 59600000.0ns 0V 59640000.0ns 0V 60440000.0ns 0V 60480000.0ns 0V 60560000.0ns 0V 60600000.0ns 0V 61400000.0ns 0V 61440000.0ns 0V 62160000.0ns 0V 62200000.0ns 0V 62680000.0ns 0V 62720000.0ns 0V 63440000.0ns 0V 63480000.0ns 0V 64280000.0ns 0V 64320000.0ns 0V 64400000.0ns 0V 64440000.0ns 0V 65240000.0ns 0V 65280000.0ns 0V 66000000.0ns 0V 66040000.0ns 0V 66520000.0ns 0V 66560000.0ns 0V 67280000.0ns 0V 67320000.0ns 0V 68120000.0ns 0V 68160000.0ns 0V 68240000.0ns 0V 68280000.0ns 0V 69080000.0ns 0V 69120000.0ns 0V 69840000.0ns 0V 69880000.0ns 0V 70360000.0ns 0V 70400000.0ns 0V 71120000.0ns 0V 71160000.0ns 0V 71960000.0ns 0V 72000000.0ns 0V 72080000.0ns 0V 72120000.0ns 0V 72920000.0ns 0V 72960000.0ns 0V 73680000.0ns 0V 73720000.0ns 0V 74200000.0ns 0V 74240000.0ns 0V 74960000.0ns 0V 75000000.0ns 0V 75800000.0ns 0V 75840000.0ns 0V 75920000.0ns 0V 75960000.0ns 0V 76760000.0ns 0V 76800000.0ns 0V 77520000.0ns 0V 77560000.0ns 0V 78040000.0ns 0V 78080000.0ns 0V 78800000.0ns 0V 78840000.0ns 0V 79640000.0ns 0V 79680000.0ns 0V 79760000.0ns 0V 79800000.0ns 0V 80600000.0ns 0V 80640000.0ns 0V 81360000.0ns 0V 81400000.0ns 0V 81880000.0ns 0V 81920000.0ns 0V 82640000.0ns 0V 82680000.0ns 0V 83480000.0ns 0V 83520000.0ns 0V 83600000.0ns 0V 83640000.0ns 0V 84440000.0ns 0V 84480000.0ns 0V 85200000.0ns 0V 85240000.0ns 0V 85720000.0ns 0V 85760000.0ns 0V 86480000.0ns 0V 86520000.0ns 0V 87320000.0ns 0V 87360000.0ns 0V 87440000.0ns 0V 87480000.0ns 0V 88280000.0ns 0V 88320000.0ns 0V 89040000.0ns 0V 89080000.0ns 0V 89560000.0ns 0V 89600000.0ns 0V 90320000.0ns 0V 90360000.0ns 0V 91160000.0ns 0V 91200000.0ns 0V 91280000.0ns 0V 91320000.0ns 0V 92120000.0ns 0V 92160000.0ns 0V 92880000.0ns 0V 92920000.0ns 0V 93400000.0ns 0V 93440000.0ns 0V 94160000.0ns 0V 94200000.0ns 0V 95000000.0ns 0V 95040000.0ns 0V 95120000.0ns 0V 95160000.0ns 0V 95960000.0ns 0V 96000000.0ns 0V 96720000.0ns 0V 96760000.0ns 0V 97240000.0ns 0V 97280000.0ns 0V 98000000.0ns 0V 98040000.0ns 0V 98840000.0ns 0V 98880000.0ns 0V 98960000.0ns 0V 99000000.0ns 0V 99800000.0ns 0V 99840000.0ns 0V 100560000.0ns 0V 100600000.0ns 0V 101080000.0ns 0V 101120000.0ns 0V 101840000.0ns 0V 101880000.0ns 0V 102680000.0ns 0V 102720000.0ns 0V 102800000.0ns 0V 102840000.0ns 0V 103640000.0ns 0V 103680000.0ns 0V 104400000.0ns 0V 104440000.0ns 0V 104920000.0ns 0V 104960000.0ns 0V 105680000.0ns 0V 105720000.0ns 0V 106520000.0ns 0V 106560000.0ns 0V 106640000.0ns 0V 106680000.0ns 0V 107480000.0ns 0V 107520000.0ns 0V 108240000.0ns 0V 108280000.0ns 0V 108760000.0ns 0V 108800000.0ns 0V 109520000.0ns 0V 109560000.0ns 0V 110360000.0ns 0V 110400000.0ns 0V 110480000.0ns 0V 110520000.0ns 0V 111320000.0ns 0V 111360000.0ns 0V 112080000.0ns 0V 112120000.0ns 0V 112600000.0ns 0V 112640000.0ns 0V 113360000.0ns 0V 113400000.0ns 0V 114200000.0ns 0V 114240000.0ns 0V 114320000.0ns 0V 114360000.0ns 0V 115160000.0ns 0V 115200000.0ns 0V 115920000.0ns 0V 115960000.0ns 0V 116440000.0ns 0V 116480000.0ns 0V 117200000.0ns 0V 117240000.0ns 0V 118040000.0ns 0V 118080000.0ns 0V 118160000.0ns 0V 118200000.0ns 0V 119000000.0ns 0V 119040000.0ns 0V 119760000.0ns 0V 119800000.0ns 0V 120280000.0ns 0V 120320000.0ns 0V 121040000.0ns 0V 121080000.0ns 0V 121880000.0ns 0V 121920000.0ns 0V 122000000.0ns 0V 122040000.0ns 0V 122840000.0ns 0V 122880000.0ns 0V 123600000.0ns 0V 123640000.0ns 0V 124120000.0ns 0V 124160000.0ns 0V 124880000.0ns 0V 124920000.0ns 0V 125720000.0ns 0V 125760000.0ns 0V 125840000.0ns 0V 125880000.0ns 0V 126680000.0ns 0V 126720000.0ns 0V 127440000.0ns 0V 127480000.0ns 0V 127960000.0ns 0V 128000000.0ns 0V 128720000.0ns 0V 128760000.0ns 0V 129560000.0ns 0V 129600000.0ns 0V 129680000.0ns 0V 129720000.0ns 0V 130520000.0ns 0V 130560000.0ns 0V 131280000.0ns 0V 131320000.0ns 0V 131800000.0ns 0V 131840000.0ns 0V 132560000.0ns 0V 132600000.0ns 0V 133400000.0ns 0V 133440000.0ns 0V 133520000.0ns 0V 133560000.0ns 0V 134360000.0ns 0V 134400000.0ns 0V 135120000.0ns 0V 135160000.0ns 0V 135640000.0ns 0V 135680000.0ns 0V 136400000.0ns 0V 136440000.0ns 0V 137240000.0ns 0V 137280000.0ns 0V 137360000.0ns 0V 137400000.0ns 0V 138200000.0ns 0V 138240000.0ns 0V 138960000.0ns 0V 139000000.0ns 0V 139480000.0ns 0V 139520000.0ns 0V 140240000.0ns 0V 140280000.0ns 0V 141080000.0ns 0V 141120000.0ns 0V 141200000.0ns 0V 141240000.0ns 0V 142040000.0ns 0V 142080000.0ns 0V 142800000.0ns 0V 142840000.0ns 0V 143320000.0ns 0V 143360000.0ns 0V 144080000.0ns 0V 144120000.0ns 0V 144920000.0ns 0V 144960000.0ns 0V 145040000.0ns 0V 145080000.0ns 0V 145880000.0ns 0V 145920000.0ns 0V 146640000.0ns 0V 146680000.0ns 0V 147160000.0ns 0V 147200000.0ns 0V 147920000.0ns 0V 147960000.0ns 0V 148760000.0ns 0V 148800000.0ns 0V 148880000.0ns 0V 148920000.0ns 0V 149720000.0ns 0V 149760000.0ns 0V 150480000.0ns 0V 150520000.0ns 0V 151000000.0ns 0V 151040000.0ns 0V 151760000.0ns 0V 151800000.0ns 0V 152600000.0ns 0V 152640000.0ns 0V 152720000.0ns 0V 152760000.0ns 0V 153560000.0ns 0V 153600000.0ns 0V 154320000.0ns 0V 154360000.0ns 0V 154840000.0ns 0V 154880000.0ns 0V 155600000.0ns 0V 155640000.0ns 0V 156440000.0ns 0V 156480000.0ns 0V 156560000.0ns 0V 156600000.0ns 0V 157400000.0ns 0V 157440000.0ns 0V 158160000.0ns 0V 158200000.0ns 0V 158680000.0ns 0V 158720000.0ns 0V 159440000.0ns 0V 159480000.0ns 0V 160280000.0ns 0V 160320000.0ns 0V 160400000.0ns 0V 160440000.0ns 0V 161240000.0ns 0V 161280000.0ns 0V 162000000.0ns 0V 162040000.0ns 0V 162520000.0ns 0V 162560000.0ns 0V 163280000.0ns 0V 163320000.0ns 0V 164120000.0ns 0V 164160000.0ns 0V 164240000.0ns 0V 164280000.0ns 0V 165080000.0ns 0V 165120000.0ns 0V 165840000.0ns 0V 165880000.0ns 0V 166360000.0ns 0V 166400000.0ns 0V 167120000.0ns 0V 167160000.0ns 0V 167960000.0ns 0V 168000000.0ns 0V 168080000.0ns 0V 168120000.0ns 0V 168920000.0ns 0V 168960000.0ns 0V 169680000.0ns 0V 169720000.0ns 0V 170200000.0ns 0V 170240000.0ns 0V 170960000.0ns 0V 171000000.0ns 0V 171800000.0ns 0V 171840000.0ns 0V 171920000.0ns 0V 171960000.0ns 0V 172760000.0ns 0V 172800000.0ns 0V 173520000.0ns 0V 173560000.0ns 0V 174040000.0ns 0V 174080000.0ns 0V 174800000.0ns 0V 174840000.0ns 0V 175640000.0ns 0V 175680000.0ns 0V 175760000.0ns 0V 175800000.0ns 0V 176600000.0ns 0V 176640000.0ns 0V 177360000.0ns 0V 177400000.0ns 0V 177880000.0ns 0V 177920000.0ns 0V 178640000.0ns 0V 178680000.0ns 0V 179480000.0ns 0V 179520000.0ns 0V 179600000.0ns 0V 179640000.0ns 0V 180440000.0ns 0V 180480000.0ns 0V 181200000.0ns 0V 181240000.0ns 0V 181720000.0ns 0V 181760000.0ns 0V 182480000.0ns 0V 182520000.0ns 0V 183320000.0ns 0V 183360000.0ns 0V 183440000.0ns 0V 183480000.0ns 0V 184280000.0ns 0V 184320000.0ns 0V 185040000.0ns 0V 185080000.0ns 0V 185560000.0ns 0V 185600000.0ns 0V 186320000.0ns 0V 186360000.0ns 0V 187160000.0ns 0V 187200000.0ns 0V 187280000.0ns 0V 187320000.0ns 0V 188120000.0ns 0V 188160000.0ns 0V 188880000.0ns 0V 188920000.0ns 0V 189400000.0ns 0V 189440000.0ns 0V 190160000.0ns 0V 190200000.0ns 0V 191000000.0ns 0V 191040000.0ns 0V 191120000.0ns 0V 191160000.0ns 0V 191960000.0ns 0V 192000000.0ns 0V 192720000.0ns 0V 192760000.0ns 0V 193240000.0ns 0V 193280000.0ns 0V 194000000.0ns 0V 194040000.0ns 0V 194840000.0ns 0V 194880000.0ns 0V 194960000.0ns 0V 195000000.0ns 0V 195800000.0ns 0V 195840000.0ns 0V 196560000.0ns 0V 196600000.0ns 0V 197080000.0ns 0V 197120000.0ns 0V 197840000.0ns 0V 197880000.0ns 0V 198680000.0ns 0V 198720000.0ns 0V 198800000.0ns 0V 198840000.0ns 0V 199640000.0ns 0V 199680000.0ns 0V 200400000.0ns 0V 200440000.0ns 0V 200920000.0ns 0V 200960000.0ns 0V 201680000.0ns 0V 201720000.0ns 0V 202520000.0ns 0V 202560000.0ns 0V 202640000.0ns 0V 202680000.0ns 0V 203480000.0ns 0V 203520000.0ns 0V 204240000.0ns 0V 204280000.0ns 0V 204760000.0ns 0V 204800000.0ns 0V 205520000.0ns 0V 205560000.0ns 0V 206360000.0ns 0V 206400000.0ns 0V 206480000.0ns 0V 206520000.0ns 0V 207320000.0ns 0V 207360000.0ns 0V 208080000.0ns 0V 208120000.0ns 0V 208600000.0ns 0V 208640000.0ns 0V 209360000.0ns 0V 209400000.0ns 0V 210200000.0ns 0V 210240000.0ns 0V 210320000.0ns 0V 210360000.0ns 0V 211160000.0ns 0V 211200000.0ns 0V 211920000.0ns 0V 211960000.0ns 0V 212440000.0ns 0V 212480000.0ns 0V 213200000.0ns 0V 213240000.0ns 0V 214040000.0ns 0V 214080000.0ns 0V 214160000.0ns 0V 214200000.0ns 0V 215000000.0ns 0V 215040000.0ns 0V 215760000.0ns 0V 215800000.0ns 0V 216280000.0ns 0V 216320000.0ns 0V 217040000.0ns 0V 217080000.0ns 0V 217880000.0ns 0V 217920000.0ns 0V 218000000.0ns 0V 218040000.0ns 0V 218840000.0ns 0V 218880000.0ns 0V 219600000.0ns 0V 219640000.0ns 0V 220120000.0ns 0V 220160000.0ns 0V 220880000.0ns 0V 220920000.0ns 0V 221720000.0ns 0V 221760000.0ns 0V 221840000.0ns 0V 221880000.0ns 0V 222680000.0ns 0V 222720000.0ns 0V 223440000.0ns 0V 223480000.0ns 0V 223960000.0ns 0V 224000000.0ns 0V 224720000.0ns 0V 224760000.0ns 0V 225560000.0ns 0V 225600000.0ns 0V 225680000.0ns 0V 225720000.0ns 0V 226520000.0ns 0V 226560000.0ns 0V 227280000.0ns 0V 227320000.0ns 0V 227800000.0ns 0V 227840000.0ns 0V 228560000.0ns 0V 228600000.0ns 0V 229400000.0ns 0V 229440000.0ns 0V 229520000.0ns 0V 229560000.0ns 0V 230360000.0ns 0V 230400000.0ns 0V 231120000.0ns 0V 231160000.0ns 0V 231640000.0ns 0V 231680000.0ns 0V 232400000.0ns 0V 232440000.0ns 0V 233240000.0ns 0V 233280000.0ns 0V 233360000.0ns 0V 233400000.0ns 0V 234200000.0ns 0V 234240000.0ns 0V 234960000.0ns 0V 235000000.0ns 0V 235480000.0ns 0V 235520000.0ns 0V 236240000.0ns 0V 236280000.0ns 0V 237080000.0ns 0V 237120000.0ns 0V 237200000.0ns 0V 237240000.0ns 0V 238040000.0ns 0V 238080000.0ns 0V 238800000.0ns 0V 238840000.0ns 0V 239320000.0ns 0V 239360000.0ns 0V 240080000.0ns 0V 240120000.0ns 0V 240920000.0ns 0V 240960000.0ns 0V 241040000.0ns 0V 241080000.0ns 0V 241880000.0ns 0V 241920000.0ns 0V 242640000.0ns 0V 242680000.0ns 0V 243160000.0ns 0V 243200000.0ns 0V 243920000.0ns 0V 243960000.0ns 0V 244760000.0ns 0V 244800000.0ns 0V 244880000.0ns 0V 244920000.0ns 0V 245720000.0ns 0V 245760000.0ns 0V 246480000.0ns 0V 246520000.0ns 0V 247000000.0ns 0V 247040000.0ns 0V 247760000.0ns 0V 247800000.0ns 0V 248600000.0ns 0V 248640000.0ns 0V 248720000.0ns 0V 248760000.0ns 0V 249560000.0ns 0V 249600000.0ns 0V 250320000.0ns 0V 250360000.0ns 0V 250840000.0ns 0V 250880000.0ns 0V 251600000.0ns 0V 251640000.0ns 0V 252440000.0ns 0V 252480000.0ns 0V 252560000.0ns 0V 252600000.0ns 0V 253400000.0ns 0V 253440000.0ns 0V 254160000.0ns 0V 254200000.0ns 0V 254680000.0ns 0V 254720000.0ns 0V 255440000.0ns 0V 255480000.0ns 0V 256280000.0ns 0V 256320000.0ns 0V 256400000.0ns 0V 256440000.0ns 0V 257240000.0ns 0V 257280000.0ns 0V 258000000.0ns 0V 258040000.0ns 0V 258520000.0ns 0V 258560000.0ns 0V 259280000.0ns 0V 259320000.0ns 0V 260120000.0ns 0V 260160000.0ns 0V 260240000.0ns 0V 260280000.0ns 0V 261080000.0ns 0V 261120000.0ns 0V 261840000.0ns 0V 261880000.0ns 0V 262360000.0ns 0V 262400000.0ns 0V 263120000.0ns 0V 263160000.0ns 0V 263960000.0ns 0V 264000000.0ns 0V 264080000.0ns 0V 264120000.0ns 0V 264920000.0ns 0V 264960000.0ns 0V 265680000.0ns 0V 265720000.0ns 0V 266200000.0ns 0V 266240000.0ns 0V 266960000.0ns 0V 267000000.0ns 0V 267800000.0ns 0V 267840000.0ns 0V 267920000.0ns 0V 267960000.0ns 0V 268760000.0ns 0V 268800000.0ns 0V 269520000.0ns 0V 269560000.0ns 0V 270040000.0ns 0V 270080000.0ns 0V 270800000.0ns 0V 270840000.0ns 0V 271640000.0ns 0V 271680000.0ns 0V 271760000.0ns 0V 271800000.0ns 0V 272600000.0ns 0V 272640000.0ns 0V 273360000.0ns 0V 273400000.0ns 0V 273880000.0ns 0V 273920000.0ns 0V 274640000.0ns 0V 274680000.0ns 0V 275480000.0ns 0V 275520000.0ns 0V 275600000.0ns 0V 275640000.0ns 0V 276440000.0ns 0V 276480000.0ns 0V 277200000.0ns 0V 277240000.0ns 0V 277720000.0ns 0V 277760000.0ns 0V 278480000.0ns 0V 278520000.0ns 0V 279320000.0ns 0V 279360000.0ns 0V 279440000.0ns 0V 279480000.0ns 0V 280280000.0ns 0V 280320000.0ns 0V 281040000.0ns 0V 281080000.0ns 0V 281560000.0ns 0V 281600000.0ns 0V 282320000.0ns 0V 282360000.0ns 0V 283160000.0ns 0V 283200000.0ns 0V 283280000.0ns 0V 283320000.0ns 0V 284120000.0ns 0V 284160000.0ns 0V 284880000.0ns 0V 284920000.0ns 0V 285400000.0ns 0V 285440000.0ns 0V 286160000.0ns 0V 286200000.0ns 0V 287000000.0ns 0V 287040000.0ns 0V 287120000.0ns 0V 287160000.0ns 0V 287960000.0ns 0V 288000000.0ns 0V 288720000.0ns 0V 288760000.0ns 0V 289240000.0ns 0V 289280000.0ns 0V 290000000.0ns 0V 290040000.0ns 0V 290840000.0ns 0V 290880000.0ns 0V 290960000.0ns 0V 291000000.0ns 0V 291800000.0ns 0V 291840000.0ns 0V 292560000.0ns 0V 292600000.0ns 0V 293080000.0ns 0V 293120000.0ns 0V 293840000.0ns 0V 293880000.0ns 0V 294680000.0ns 0V 294720000.0ns 0V 294800000.0ns 0V 294840000.0ns 0V 295640000.0ns 0V 295680000.0ns 0V 296400000.0ns 0V 296440000.0ns 0V 296920000.0ns 0V 296960000.0ns 0V 297680000.0ns 0V 297720000.0ns 0V 298520000.0ns 0V 298560000.0ns 0V 298640000.0ns 0V 298680000.0ns 0V 299480000.0ns 0V 299520000.0ns 0V 300240000.0ns 0V 300280000.0ns 0V 300760000.0ns 0V 300800000.0ns 0V 301520000.0ns 0V 301560000.0ns 0V 302360000.0ns 0V 302400000.0ns 0V 302480000.0ns 0V 302520000.0ns 0V 303320000.0ns 0V 303360000.0ns 0V 304080000.0ns 0V 304120000.0ns 0V 304600000.0ns 0V 304640000.0ns 0V 305360000.0ns 0V 305400000.0ns 0V 306200000.0ns 0V 306240000.0ns 0V 306320000.0ns 0V 306360000.0ns 0V 307160000.0ns 0V 307200000.0ns 0V 307920000.0ns 0V 307960000.0ns 0V 308440000.0ns 0V 308480000.0ns 0V 309200000.0ns 0V 309240000.0ns 0V 310040000.0ns 0V 310080000.0ns 0V 310160000.0ns 0V 310200000.0ns 0V 311000000.0ns 0V 311040000.0ns 0V 311760000.0ns 0V 311800000.0ns 0V 312280000.0ns 0V 312320000.0ns 0V 313040000.0ns 0V 313080000.0ns 0V 313880000.0ns 0V 313920000.0ns 0V 314000000.0ns 0V 314040000.0ns 0V 314840000.0ns 0V 314880000.0ns 0V 315600000.0ns 0V 315640000.0ns 0V 316120000.0ns 0V 316160000.0ns 0V 316880000.0ns 0V 316920000.0ns 0V 317720000.0ns 0V 317760000.0ns 0V 317840000.0ns 0V 317880000.0ns 0V 318680000.0ns 0V 318720000.0ns 0V 319440000.0ns 0V 319480000.0ns 0V 319960000.0ns 0V 320000000.0ns 0V 320720000.0ns 0V 320760000.0ns 0V 321560000.0ns 0V 321600000.0ns 0V 321680000.0ns 0V 321720000.0ns 0V 322520000.0ns 0V 322560000.0ns 0V 323280000.0ns 0V 323320000.0ns 0V 323800000.0ns 0V 323840000.0ns 0V 324560000.0ns 0V 324600000.0ns 0V 325400000.0ns 0V 325440000.0ns 0V 325520000.0ns 0V 325560000.0ns 0V 326360000.0ns 0V 326400000.0ns 0V 327120000.0ns 0V 327160000.0ns 0V 327640000.0ns 0V 327680000.0ns 0V 328400000.0ns 0V 328440000.0ns 0V 329240000.0ns 0V 329280000.0ns 0V 329360000.0ns 0V 329400000.0ns 0V 330200000.0ns 0V 330240000.0ns 0V 330960000.0ns 0V 331000000.0ns 0V 331480000.0ns 0V 331520000.0ns 0V 332240000.0ns 0V 332280000.0ns 0V 333080000.0ns 0V 333120000.0ns 0V 333200000.0ns 0V 333240000.0ns 0V 334040000.0ns 0V 334080000.0ns 0V 334800000.0ns 0V 334840000.0ns 0V 335320000.0ns 0V 335360000.0ns 0V 336080000.0ns 0V 336120000.0ns 0V 336920000.0ns 0V 336960000.0ns 0V 337040000.0ns 0V 337080000.0ns 0V 337880000.0ns 0V 337920000.0ns 0V 338640000.0ns 0V 338680000.0ns 0V 339160000.0ns 0V 339200000.0ns 0V 339920000.0ns 0V 339960000.0ns 0V 340760000.0ns 0V 340800000.0ns 0V 340880000.0ns 0V 340920000.0ns 0V 341720000.0ns 0V 341760000.0ns 0V 342480000.0ns 0V 342520000.0ns 0V 343000000.0ns 0V 343040000.0ns 0V 343760000.0ns 0V 343800000.0ns 0V 344600000.0ns 0V 344640000.0ns 0V 344720000.0ns 0V 344760000.0ns 0V 345560000.0ns 0V 345600000.0ns 0V 346320000.0ns 0V 346360000.0ns 0V 346840000.0ns 0V 346880000.0ns 0V 347600000.0ns 0V 347640000.0ns 0V 348440000.0ns 0V 348480000.0ns 0V 348560000.0ns 0V 348600000.0ns 0V 349400000.0ns 0V 349440000.0ns 0V 350160000.0ns 0V 350200000.0ns 0V 350680000.0ns 0V 350720000.0ns 0V 351440000.0ns 0V 351480000.0ns 0V 352280000.0ns 0V 352320000.0ns 0V 352400000.0ns 0V 352440000.0ns 0V 353240000.0ns 0V 353280000.0ns 0V 354000000.0ns 0V 354040000.0ns 0V 354520000.0ns 0V 354560000.0ns 0V 355280000.0ns 0V 355320000.0ns 0V 356120000.0ns 0V 356160000.0ns 0V 356240000.0ns 0V 356280000.0ns 0V 357080000.0ns 0V 357120000.0ns 0V 357840000.0ns 0V 357880000.0ns 0V 358360000.0ns 0V 358400000.0ns 0V 359120000.0ns 0V 359160000.0ns 0V 359960000.0ns 0V 360000000.0ns 0V 360080000.0ns 0V 360120000.0ns 0V 360920000.0ns 0V 360960000.0ns 0V 361680000.0ns 0V 361720000.0ns 0V 362200000.0ns 0V 362240000.0ns 0V 362960000.0ns 0V 363000000.0ns 0V 363800000.0ns 0V 363840000.0ns 0V 363920000.0ns 0V 363960000.0ns 0V 364760000.0ns 0V 364800000.0ns 0V 365520000.0ns 0V 365560000.0ns 0V 366040000.0ns 0V 366080000.0ns 0V 366800000.0ns 0V 366840000.0ns 0V 367640000.0ns 0V 367680000.0ns 0V 367760000.0ns 0V 367800000.0ns 0V 368600000.0ns 0V 368640000.0ns 0V 369360000.0ns 0V 369400000.0ns 0V 369880000.0ns 0V 369920000.0ns 0V 370640000.0ns 0V 370680000.0ns 0V 371480000.0ns 0V 371520000.0ns 0V 371600000.0ns 0V 371640000.0ns 0V 372440000.0ns 0V 372480000.0ns 0V 373200000.0ns 0V 373240000.0ns 0V 373720000.0ns 0V 373760000.0ns 0V 374480000.0ns 0V 374520000.0ns 0V 375320000.0ns 0V 375360000.0ns 0V 375440000.0ns 0V 375480000.0ns 0V 376280000.0ns 0V 376320000.0ns 0V 377040000.0ns 0V 377080000.0ns 0V 377560000.0ns 0V 377600000.0ns 0V 378320000.0ns 0V 378360000.0ns 0V 379160000.0ns 0V 379200000.0ns 0V 379280000.0ns 0V 379320000.0ns 0V 380120000.0ns 0V 380160000.0ns 0V 380880000.0ns 0V 380920000.0ns 0V 381400000.0ns 0V 381440000.0ns 0V 382160000.0ns 0V 382200000.0ns 0V 383000000.0ns 0V 383040000.0ns 0V 383120000.0ns 0V 383160000.0ns 0V 383960000.0ns 0V 384000000.0ns 0V 384720000.0ns 0V 384760000.0ns 0V 385240000.0ns 0V 385280000.0ns 0V 386000000.0ns 0V 386040000.0ns 0V 386840000.0ns 0V 386880000.0ns 0V 386960000.0ns 0V 387000000.0ns 0V 387800000.0ns 0V 387840000.0ns 0V 388560000.0ns 0V 388600000.0ns 0V 389080000.0ns 0V 389120000.0ns 0V 389840000.0ns 0V 389880000.0ns 0V 390680000.0ns 0V 390720000.0ns 0V 390800000.0ns 0V 390840000.0ns 0V)
VVWWL_I2 WWL_I2 0 PWL(0ns 0V 1800000.0ns 0V 1840000.0ns 1.95V 2240000.0ns 1.95V 2280000.0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0V 8400000.0ns 0V 8440000.0ns 0V 8920000.0ns 0V 8960000.0ns 0V 9680000.0ns 0V 9720000.0ns 0V 10520000.0ns 0V 10560000.0ns 0V 10640000.0ns 0V 10680000.0ns 0V 11480000.0ns 0V 11520000.0ns 0V 12240000.0ns 0V 12280000.0ns 0V 12760000.0ns 0V 12800000.0ns 0V 13520000.0ns 0V 13560000.0ns 0V 14360000.0ns 0V 14400000.0ns 0V 14480000.0ns 0V 14520000.0ns 0V 15320000.0ns 0V 15360000.0ns 0V 16080000.0ns 0V 16120000.0ns 0V 16600000.0ns 0V 16640000.0ns 0V 17360000.0ns 0V 17400000.0ns 0V 18200000.0ns 0V 18240000.0ns 0V 18320000.0ns 0V 18360000.0ns 0V 19160000.0ns 0V 19200000.0ns 0V 19920000.0ns 0V 19960000.0ns 0V 20440000.0ns 0V 20480000.0ns 0V 21200000.0ns 0V 21240000.0ns 0V 22040000.0ns 0V 22080000.0ns 0V 22160000.0ns 0V 22200000.0ns 0V 23000000.0ns 0V 23040000.0ns 0V 23760000.0ns 0V 23800000.0ns 0V 24280000.0ns 0V 24320000.0ns 0V 25040000.0ns 0V 25080000.0ns 0V 25880000.0ns 0V 25920000.0ns 0V 26000000.0ns 0V 26040000.0ns 0V 26840000.0ns 0V 26880000.0ns 0V 27600000.0ns 0V 27640000.0ns 0V 28120000.0ns 0V 28160000.0ns 0V 28880000.0ns 0V 28920000.0ns 0V 29720000.0ns 0V 29760000.0ns 0V 29840000.0ns 0V 29880000.0ns 0V 30680000.0ns 0V 30720000.0ns 0V 31440000.0ns 0V 31480000.0ns 0V 31960000.0ns 0V 32000000.0ns 0V 32720000.0ns 0V 32760000.0ns 0V 33560000.0ns 0V 33600000.0ns 0V 33680000.0ns 0V 33720000.0ns 0V 34520000.0ns 0V 34560000.0ns 0V 35280000.0ns 0V 35320000.0ns 0V 35800000.0ns 0V 35840000.0ns 0V 36560000.0ns 0V 36600000.0ns 0V 37400000.0ns 0V 37440000.0ns 0V 37520000.0ns 0V 37560000.0ns 0V 38360000.0ns 0V 38400000.0ns 0V 39120000.0ns 0V 39160000.0ns 0V 39640000.0ns 0V 39680000.0ns 0V 40400000.0ns 0V 40440000.0ns 0V 41240000.0ns 0V 41280000.0ns 0V 41360000.0ns 0V 41400000.0ns 0V 42200000.0ns 0V 42240000.0ns 0V 42960000.0ns 0V 43000000.0ns 0V 43480000.0ns 0V 43520000.0ns 0V 44240000.0ns 0V 44280000.0ns 0V 45080000.0ns 0V 45120000.0ns 0V 45200000.0ns 0V 45240000.0ns 0V 46040000.0ns 0V 46080000.0ns 0V 46800000.0ns 0V 46840000.0ns 0V 47320000.0ns 0V 47360000.0ns 0V 48080000.0ns 0V 48120000.0ns 0V 48920000.0ns 0V 48960000.0ns 0V 49040000.0ns 0V 49080000.0ns 0V 49880000.0ns 0V 49920000.0ns 0V 50640000.0ns 0V 50680000.0ns 0V 51160000.0ns 0V 51200000.0ns 0V 51920000.0ns 0V 51960000.0ns 0V 52760000.0ns 0V 52800000.0ns 0V 52880000.0ns 0V 52920000.0ns 0V 53720000.0ns 0V 53760000.0ns 0V 54480000.0ns 0V 54520000.0ns 0V 55000000.0ns 0V 55040000.0ns 0V 55760000.0ns 0V 55800000.0ns 0V 56600000.0ns 0V 56640000.0ns 0V 56720000.0ns 0V 56760000.0ns 0V 57560000.0ns 0V 57600000.0ns 0V 58320000.0ns 0V 58360000.0ns 0V 58840000.0ns 0V 58880000.0ns 0V 59600000.0ns 0V 59640000.0ns 0V 60440000.0ns 0V 60480000.0ns 0V 60560000.0ns 0V 60600000.0ns 0V 61400000.0ns 0V 61440000.0ns 0V 62160000.0ns 0V 62200000.0ns 0V 62680000.0ns 0V 62720000.0ns 0V 63440000.0ns 0V 63480000.0ns 0V 64280000.0ns 0V 64320000.0ns 0V 64400000.0ns 0V 64440000.0ns 0V 65240000.0ns 0V 65280000.0ns 0V 66000000.0ns 0V 66040000.0ns 0V 66520000.0ns 0V 66560000.0ns 0V 67280000.0ns 0V 67320000.0ns 0V 68120000.0ns 0V 68160000.0ns 0V 68240000.0ns 0V 68280000.0ns 0V 69080000.0ns 0V 69120000.0ns 0V 69840000.0ns 0V 69880000.0ns 0V 70360000.0ns 0V 70400000.0ns 0V 71120000.0ns 0V 71160000.0ns 0V 71960000.0ns 0V 72000000.0ns 0V 72080000.0ns 0V 72120000.0ns 0V 72920000.0ns 0V 72960000.0ns 0V 73680000.0ns 0V 73720000.0ns 0V 74200000.0ns 0V 74240000.0ns 0V 74960000.0ns 0V 75000000.0ns 0V 75800000.0ns 0V 75840000.0ns 0V 75920000.0ns 0V 75960000.0ns 0V 76760000.0ns 0V 76800000.0ns 0V 77520000.0ns 0V 77560000.0ns 0V 78040000.0ns 0V 78080000.0ns 0V 78800000.0ns 0V 78840000.0ns 0V 79640000.0ns 0V 79680000.0ns 0V 79760000.0ns 0V 79800000.0ns 0V 80600000.0ns 0V 80640000.0ns 0V 81360000.0ns 0V 81400000.0ns 0V 81880000.0ns 0V 81920000.0ns 0V 82640000.0ns 0V 82680000.0ns 0V 83480000.0ns 0V 83520000.0ns 0V 83600000.0ns 0V 83640000.0ns 0V 84440000.0ns 0V 84480000.0ns 0V 85200000.0ns 0V 85240000.0ns 0V 85720000.0ns 0V 85760000.0ns 0V 86480000.0ns 0V 86520000.0ns 0V 87320000.0ns 0V 87360000.0ns 0V 87440000.0ns 0V 87480000.0ns 0V 88280000.0ns 0V 88320000.0ns 0V 89040000.0ns 0V 89080000.0ns 0V 89560000.0ns 0V 89600000.0ns 0V 90320000.0ns 0V 90360000.0ns 0V 91160000.0ns 0V 91200000.0ns 0V 91280000.0ns 0V 91320000.0ns 0V 92120000.0ns 0V 92160000.0ns 0V 92880000.0ns 0V 92920000.0ns 0V 93400000.0ns 0V 93440000.0ns 0V 94160000.0ns 0V 94200000.0ns 0V 95000000.0ns 0V 95040000.0ns 0V 95120000.0ns 0V 95160000.0ns 0V 95960000.0ns 0V 96000000.0ns 0V 96720000.0ns 0V 96760000.0ns 0V 97240000.0ns 0V 97280000.0ns 0V 98000000.0ns 0V 98040000.0ns 0V 98840000.0ns 0V 98880000.0ns 0V 98960000.0ns 0V 99000000.0ns 0V 99800000.0ns 0V 99840000.0ns 0V 100560000.0ns 0V 100600000.0ns 0V 101080000.0ns 0V 101120000.0ns 0V 101840000.0ns 0V 101880000.0ns 0V 102680000.0ns 0V 102720000.0ns 0V 102800000.0ns 0V 102840000.0ns 0V 103640000.0ns 0V 103680000.0ns 0V 104400000.0ns 0V 104440000.0ns 0V 104920000.0ns 0V 104960000.0ns 0V 105680000.0ns 0V 105720000.0ns 0V 106520000.0ns 0V 106560000.0ns 0V 106640000.0ns 0V 106680000.0ns 0V 107480000.0ns 0V 107520000.0ns 0V 108240000.0ns 0V 108280000.0ns 0V 108760000.0ns 0V 108800000.0ns 0V 109520000.0ns 0V 109560000.0ns 0V 110360000.0ns 0V 110400000.0ns 0V 110480000.0ns 0V 110520000.0ns 0V 111320000.0ns 0V 111360000.0ns 0V 112080000.0ns 0V 112120000.0ns 0V 112600000.0ns 0V 112640000.0ns 0V 113360000.0ns 0V 113400000.0ns 0V 114200000.0ns 0V 114240000.0ns 0V 114320000.0ns 0V 114360000.0ns 0V 115160000.0ns 0V 115200000.0ns 0V 115920000.0ns 0V 115960000.0ns 0V 116440000.0ns 0V 116480000.0ns 0V 117200000.0ns 0V 117240000.0ns 0V 118040000.0ns 0V 118080000.0ns 0V 118160000.0ns 0V 118200000.0ns 0V 119000000.0ns 0V 119040000.0ns 0V 119760000.0ns 0V 119800000.0ns 0V 120280000.0ns 0V 120320000.0ns 0V 121040000.0ns 0V 121080000.0ns 0V 121880000.0ns 0V 121920000.0ns 0V 122000000.0ns 0V 122040000.0ns 0V 122840000.0ns 0V 122880000.0ns 0V 123600000.0ns 0V 123640000.0ns 0V 124120000.0ns 0V 124160000.0ns 0V 124880000.0ns 0V 124920000.0ns 0V 125720000.0ns 0V 125760000.0ns 0V 125840000.0ns 0V 125880000.0ns 0V 126680000.0ns 0V 126720000.0ns 0V 127440000.0ns 0V 127480000.0ns 0V 127960000.0ns 0V 128000000.0ns 0V 128720000.0ns 0V 128760000.0ns 0V 129560000.0ns 0V 129600000.0ns 0V 129680000.0ns 0V 129720000.0ns 0V 130520000.0ns 0V 130560000.0ns 0V 131280000.0ns 0V 131320000.0ns 0V 131800000.0ns 0V 131840000.0ns 0V 132560000.0ns 0V 132600000.0ns 0V 133400000.0ns 0V 133440000.0ns 0V 133520000.0ns 0V 133560000.0ns 0V 134360000.0ns 0V 134400000.0ns 0V 135120000.0ns 0V 135160000.0ns 0V 135640000.0ns 0V 135680000.0ns 0V 136400000.0ns 0V 136440000.0ns 0V 137240000.0ns 0V 137280000.0ns 0V 137360000.0ns 0V 137400000.0ns 0V 138200000.0ns 0V 138240000.0ns 0V 138960000.0ns 0V 139000000.0ns 0V 139480000.0ns 0V 139520000.0ns 0V 140240000.0ns 0V 140280000.0ns 0V 141080000.0ns 0V 141120000.0ns 0V 141200000.0ns 0V 141240000.0ns 0V 142040000.0ns 0V 142080000.0ns 0V 142800000.0ns 0V 142840000.0ns 0V 143320000.0ns 0V 143360000.0ns 0V 144080000.0ns 0V 144120000.0ns 0V 144920000.0ns 0V 144960000.0ns 0V 145040000.0ns 0V 145080000.0ns 0V 145880000.0ns 0V 145920000.0ns 0V 146640000.0ns 0V 146680000.0ns 0V 147160000.0ns 0V 147200000.0ns 0V 147920000.0ns 0V 147960000.0ns 0V 148760000.0ns 0V 148800000.0ns 0V 148880000.0ns 0V 148920000.0ns 0V 149720000.0ns 0V 149760000.0ns 0V 150480000.0ns 0V 150520000.0ns 0V 151000000.0ns 0V 151040000.0ns 0V 151760000.0ns 0V 151800000.0ns 0V 152600000.0ns 0V 152640000.0ns 0V 152720000.0ns 0V 152760000.0ns 0V 153560000.0ns 0V 153600000.0ns 0V 154320000.0ns 0V 154360000.0ns 0V 154840000.0ns 0V 154880000.0ns 0V 155600000.0ns 0V 155640000.0ns 0V 156440000.0ns 0V 156480000.0ns 0V 156560000.0ns 0V 156600000.0ns 0V 157400000.0ns 0V 157440000.0ns 0V 158160000.0ns 0V 158200000.0ns 0V 158680000.0ns 0V 158720000.0ns 0V 159440000.0ns 0V 159480000.0ns 0V 160280000.0ns 0V 160320000.0ns 0V 160400000.0ns 0V 160440000.0ns 0V 161240000.0ns 0V 161280000.0ns 0V 162000000.0ns 0V 162040000.0ns 0V 162520000.0ns 0V 162560000.0ns 0V 163280000.0ns 0V 163320000.0ns 0V 164120000.0ns 0V 164160000.0ns 0V 164240000.0ns 0V 164280000.0ns 0V 165080000.0ns 0V 165120000.0ns 0V 165840000.0ns 0V 165880000.0ns 0V 166360000.0ns 0V 166400000.0ns 0V 167120000.0ns 0V 167160000.0ns 0V 167960000.0ns 0V 168000000.0ns 0V 168080000.0ns 0V 168120000.0ns 0V 168920000.0ns 0V 168960000.0ns 0V 169680000.0ns 0V 169720000.0ns 0V 170200000.0ns 0V 170240000.0ns 0V 170960000.0ns 0V 171000000.0ns 0V 171800000.0ns 0V 171840000.0ns 0V 171920000.0ns 0V 171960000.0ns 0V 172760000.0ns 0V 172800000.0ns 0V 173520000.0ns 0V 173560000.0ns 0V 174040000.0ns 0V 174080000.0ns 0V 174800000.0ns 0V 174840000.0ns 0V 175640000.0ns 0V 175680000.0ns 0V 175760000.0ns 0V 175800000.0ns 0V 176600000.0ns 0V 176640000.0ns 0V 177360000.0ns 0V 177400000.0ns 0V 177880000.0ns 0V 177920000.0ns 0V 178640000.0ns 0V 178680000.0ns 0V 179480000.0ns 0V 179520000.0ns 0V 179600000.0ns 0V 179640000.0ns 0V 180440000.0ns 0V 180480000.0ns 0V 181200000.0ns 0V 181240000.0ns 0V 181720000.0ns 0V 181760000.0ns 0V 182480000.0ns 0V 182520000.0ns 0V 183320000.0ns 0V 183360000.0ns 0V 183440000.0ns 0V 183480000.0ns 0V 184280000.0ns 0V 184320000.0ns 0V 185040000.0ns 0V 185080000.0ns 0V 185560000.0ns 0V 185600000.0ns 0V 186320000.0ns 0V 186360000.0ns 0V 187160000.0ns 0V 187200000.0ns 0V 187280000.0ns 0V 187320000.0ns 0V 188120000.0ns 0V 188160000.0ns 0V 188880000.0ns 0V 188920000.0ns 0V 189400000.0ns 0V 189440000.0ns 0V 190160000.0ns 0V 190200000.0ns 0V 191000000.0ns 0V 191040000.0ns 0V 191120000.0ns 0V 191160000.0ns 0V 191960000.0ns 0V 192000000.0ns 0V 192720000.0ns 0V 192760000.0ns 0V 193240000.0ns 0V 193280000.0ns 0V 194000000.0ns 0V 194040000.0ns 0V 194840000.0ns 0V 194880000.0ns 0V 194960000.0ns 0V 195000000.0ns 0V 195800000.0ns 0V 195840000.0ns 0V 196560000.0ns 0V 196600000.0ns 0V 197080000.0ns 0V 197120000.0ns 0V 197840000.0ns 0V 197880000.0ns 0V 198680000.0ns 0V 198720000.0ns 0V 198800000.0ns 0V 198840000.0ns 0V 199640000.0ns 0V 199680000.0ns 0V 200400000.0ns 0V 200440000.0ns 0V 200920000.0ns 0V 200960000.0ns 0V 201680000.0ns 0V 201720000.0ns 0V 202520000.0ns 0V 202560000.0ns 0V 202640000.0ns 0V 202680000.0ns 0V 203480000.0ns 0V 203520000.0ns 0V 204240000.0ns 0V 204280000.0ns 0V 204760000.0ns 0V 204800000.0ns 0V 205520000.0ns 0V 205560000.0ns 0V 206360000.0ns 0V 206400000.0ns 0V 206480000.0ns 0V 206520000.0ns 0V 207320000.0ns 0V 207360000.0ns 0V 208080000.0ns 0V 208120000.0ns 0V 208600000.0ns 0V 208640000.0ns 0V 209360000.0ns 0V 209400000.0ns 0V 210200000.0ns 0V 210240000.0ns 0V 210320000.0ns 0V 210360000.0ns 0V 211160000.0ns 0V 211200000.0ns 0V 211920000.0ns 0V 211960000.0ns 0V 212440000.0ns 0V 212480000.0ns 0V 213200000.0ns 0V 213240000.0ns 0V 214040000.0ns 0V 214080000.0ns 0V 214160000.0ns 0V 214200000.0ns 0V 215000000.0ns 0V 215040000.0ns 0V 215760000.0ns 0V 215800000.0ns 0V 216280000.0ns 0V 216320000.0ns 0V 217040000.0ns 0V 217080000.0ns 0V 217880000.0ns 0V 217920000.0ns 0V 218000000.0ns 0V 218040000.0ns 0V 218840000.0ns 0V 218880000.0ns 0V 219600000.0ns 0V 219640000.0ns 0V 220120000.0ns 0V 220160000.0ns 0V 220880000.0ns 0V 220920000.0ns 0V 221720000.0ns 0V 221760000.0ns 0V 221840000.0ns 0V 221880000.0ns 0V 222680000.0ns 0V 222720000.0ns 0V 223440000.0ns 0V 223480000.0ns 0V 223960000.0ns 0V 224000000.0ns 0V 224720000.0ns 0V 224760000.0ns 0V 225560000.0ns 0V 225600000.0ns 0V 225680000.0ns 0V 225720000.0ns 0V 226520000.0ns 0V 226560000.0ns 0V 227280000.0ns 0V 227320000.0ns 0V 227800000.0ns 0V 227840000.0ns 0V 228560000.0ns 0V 228600000.0ns 0V 229400000.0ns 0V 229440000.0ns 0V 229520000.0ns 0V 229560000.0ns 0V 230360000.0ns 0V 230400000.0ns 0V 231120000.0ns 0V 231160000.0ns 0V 231640000.0ns 0V 231680000.0ns 0V 232400000.0ns 0V 232440000.0ns 0V 233240000.0ns 0V 233280000.0ns 0V 233360000.0ns 0V 233400000.0ns 0V 234200000.0ns 0V 234240000.0ns 0V 234960000.0ns 0V 235000000.0ns 0V 235480000.0ns 0V 235520000.0ns 0V 236240000.0ns 0V 236280000.0ns 0V 237080000.0ns 0V 237120000.0ns 0V 237200000.0ns 0V 237240000.0ns 0V 238040000.0ns 0V 238080000.0ns 0V 238800000.0ns 0V 238840000.0ns 0V 239320000.0ns 0V 239360000.0ns 0V 240080000.0ns 0V 240120000.0ns 0V 240920000.0ns 0V 240960000.0ns 0V 241040000.0ns 0V 241080000.0ns 0V 241880000.0ns 0V 241920000.0ns 0V 242640000.0ns 0V 242680000.0ns 0V 243160000.0ns 0V 243200000.0ns 0V 243920000.0ns 0V 243960000.0ns 0V 244760000.0ns 0V 244800000.0ns 0V 244880000.0ns 0V 244920000.0ns 0V 245720000.0ns 0V 245760000.0ns 0V 246480000.0ns 0V 246520000.0ns 0V 247000000.0ns 0V 247040000.0ns 0V 247760000.0ns 0V 247800000.0ns 0V 248600000.0ns 0V 248640000.0ns 0V 248720000.0ns 0V 248760000.0ns 0V 249560000.0ns 0V 249600000.0ns 0V 250320000.0ns 0V 250360000.0ns 0V 250840000.0ns 0V 250880000.0ns 0V 251600000.0ns 0V 251640000.0ns 0V 252440000.0ns 0V 252480000.0ns 0V 252560000.0ns 0V 252600000.0ns 0V 253400000.0ns 0V 253440000.0ns 0V 254160000.0ns 0V 254200000.0ns 0V 254680000.0ns 0V 254720000.0ns 0V 255440000.0ns 0V 255480000.0ns 0V 256280000.0ns 0V 256320000.0ns 0V 256400000.0ns 0V 256440000.0ns 0V 257240000.0ns 0V 257280000.0ns 0V 258000000.0ns 0V 258040000.0ns 0V 258520000.0ns 0V 258560000.0ns 0V 259280000.0ns 0V 259320000.0ns 0V 260120000.0ns 0V 260160000.0ns 0V 260240000.0ns 0V 260280000.0ns 0V 261080000.0ns 0V 261120000.0ns 0V 261840000.0ns 0V 261880000.0ns 0V 262360000.0ns 0V 262400000.0ns 0V 263120000.0ns 0V 263160000.0ns 0V 263960000.0ns 0V 264000000.0ns 0V 264080000.0ns 0V 264120000.0ns 0V 264920000.0ns 0V 264960000.0ns 0V 265680000.0ns 0V 265720000.0ns 0V 266200000.0ns 0V 266240000.0ns 0V 266960000.0ns 0V 267000000.0ns 0V 267800000.0ns 0V 267840000.0ns 0V 267920000.0ns 0V 267960000.0ns 0V 268760000.0ns 0V 268800000.0ns 0V 269520000.0ns 0V 269560000.0ns 0V 270040000.0ns 0V 270080000.0ns 0V 270800000.0ns 0V 270840000.0ns 0V 271640000.0ns 0V 271680000.0ns 0V 271760000.0ns 0V 271800000.0ns 0V 272600000.0ns 0V 272640000.0ns 0V 273360000.0ns 0V 273400000.0ns 0V 273880000.0ns 0V 273920000.0ns 0V 274640000.0ns 0V 274680000.0ns 0V 275480000.0ns 0V 275520000.0ns 0V 275600000.0ns 0V 275640000.0ns 0V 276440000.0ns 0V 276480000.0ns 0V 277200000.0ns 0V 277240000.0ns 0V 277720000.0ns 0V 277760000.0ns 0V 278480000.0ns 0V 278520000.0ns 0V 279320000.0ns 0V 279360000.0ns 0V 279440000.0ns 0V 279480000.0ns 0V 280280000.0ns 0V 280320000.0ns 0V 281040000.0ns 0V 281080000.0ns 0V 281560000.0ns 0V 281600000.0ns 0V 282320000.0ns 0V 282360000.0ns 0V 283160000.0ns 0V 283200000.0ns 0V 283280000.0ns 0V 283320000.0ns 0V 284120000.0ns 0V 284160000.0ns 0V 284880000.0ns 0V 284920000.0ns 0V 285400000.0ns 0V 285440000.0ns 0V 286160000.0ns 0V 286200000.0ns 0V 287000000.0ns 0V 287040000.0ns 0V 287120000.0ns 0V 287160000.0ns 0V 287960000.0ns 0V 288000000.0ns 0V 288720000.0ns 0V 288760000.0ns 0V 289240000.0ns 0V 289280000.0ns 0V 290000000.0ns 0V 290040000.0ns 0V 290840000.0ns 0V 290880000.0ns 0V 290960000.0ns 0V 291000000.0ns 0V 291800000.0ns 0V 291840000.0ns 0V 292560000.0ns 0V 292600000.0ns 0V 293080000.0ns 0V 293120000.0ns 0V 293840000.0ns 0V 293880000.0ns 0V 294680000.0ns 0V 294720000.0ns 0V 294800000.0ns 0V 294840000.0ns 0V 295640000.0ns 0V 295680000.0ns 0V 296400000.0ns 0V 296440000.0ns 0V 296920000.0ns 0V 296960000.0ns 0V 297680000.0ns 0V 297720000.0ns 0V 298520000.0ns 0V 298560000.0ns 0V 298640000.0ns 0V 298680000.0ns 0V 299480000.0ns 0V 299520000.0ns 0V 300240000.0ns 0V 300280000.0ns 0V 300760000.0ns 0V 300800000.0ns 0V 301520000.0ns 0V 301560000.0ns 0V 302360000.0ns 0V 302400000.0ns 0V 302480000.0ns 0V 302520000.0ns 0V 303320000.0ns 0V 303360000.0ns 0V 304080000.0ns 0V 304120000.0ns 0V 304600000.0ns 0V 304640000.0ns 0V 305360000.0ns 0V 305400000.0ns 0V 306200000.0ns 0V 306240000.0ns 0V 306320000.0ns 0V 306360000.0ns 0V 307160000.0ns 0V 307200000.0ns 0V 307920000.0ns 0V 307960000.0ns 0V 308440000.0ns 0V 308480000.0ns 0V 309200000.0ns 0V 309240000.0ns 0V 310040000.0ns 0V 310080000.0ns 0V 310160000.0ns 0V 310200000.0ns 0V 311000000.0ns 0V 311040000.0ns 0V 311760000.0ns 0V 311800000.0ns 0V 312280000.0ns 0V 312320000.0ns 0V 313040000.0ns 0V 313080000.0ns 0V 313880000.0ns 0V 313920000.0ns 0V 314000000.0ns 0V 314040000.0ns 0V 314840000.0ns 0V 314880000.0ns 0V 315600000.0ns 0V 315640000.0ns 0V 316120000.0ns 0V 316160000.0ns 0V 316880000.0ns 0V 316920000.0ns 0V 317720000.0ns 0V 317760000.0ns 0V 317840000.0ns 0V 317880000.0ns 0V 318680000.0ns 0V 318720000.0ns 0V 319440000.0ns 0V 319480000.0ns 0V 319960000.0ns 0V 320000000.0ns 0V 320720000.0ns 0V 320760000.0ns 0V 321560000.0ns 0V 321600000.0ns 0V 321680000.0ns 0V 321720000.0ns 0V 322520000.0ns 0V 322560000.0ns 0V 323280000.0ns 0V 323320000.0ns 0V 323800000.0ns 0V 323840000.0ns 0V 324560000.0ns 0V 324600000.0ns 0V 325400000.0ns 0V 325440000.0ns 0V 325520000.0ns 0V 325560000.0ns 0V 326360000.0ns 0V 326400000.0ns 0V 327120000.0ns 0V 327160000.0ns 0V 327640000.0ns 0V 327680000.0ns 0V 328400000.0ns 0V 328440000.0ns 0V 329240000.0ns 0V 329280000.0ns 0V 329360000.0ns 0V 329400000.0ns 0V 330200000.0ns 0V 330240000.0ns 0V 330960000.0ns 0V 331000000.0ns 0V 331480000.0ns 0V 331520000.0ns 0V 332240000.0ns 0V 332280000.0ns 0V 333080000.0ns 0V 333120000.0ns 0V 333200000.0ns 0V 333240000.0ns 0V 334040000.0ns 0V 334080000.0ns 0V 334800000.0ns 0V 334840000.0ns 0V 335320000.0ns 0V 335360000.0ns 0V 336080000.0ns 0V 336120000.0ns 0V 336920000.0ns 0V 336960000.0ns 0V 337040000.0ns 0V 337080000.0ns 0V 337880000.0ns 0V 337920000.0ns 0V 338640000.0ns 0V 338680000.0ns 0V 339160000.0ns 0V 339200000.0ns 0V 339920000.0ns 0V 339960000.0ns 0V 340760000.0ns 0V 340800000.0ns 0V 340880000.0ns 0V 340920000.0ns 0V 341720000.0ns 0V 341760000.0ns 0V 342480000.0ns 0V 342520000.0ns 0V 343000000.0ns 0V 343040000.0ns 0V 343760000.0ns 0V 343800000.0ns 0V 344600000.0ns 0V 344640000.0ns 0V 344720000.0ns 0V 344760000.0ns 0V 345560000.0ns 0V 345600000.0ns 0V 346320000.0ns 0V 346360000.0ns 0V 346840000.0ns 0V 346880000.0ns 0V 347600000.0ns 0V 347640000.0ns 0V 348440000.0ns 0V 348480000.0ns 0V 348560000.0ns 0V 348600000.0ns 0V 349400000.0ns 0V 349440000.0ns 0V 350160000.0ns 0V 350200000.0ns 0V 350680000.0ns 0V 350720000.0ns 0V 351440000.0ns 0V 351480000.0ns 0V 352280000.0ns 0V 352320000.0ns 0V 352400000.0ns 0V 352440000.0ns 0V 353240000.0ns 0V 353280000.0ns 0V 354000000.0ns 0V 354040000.0ns 0V 354520000.0ns 0V 354560000.0ns 0V 355280000.0ns 0V 355320000.0ns 0V 356120000.0ns 0V 356160000.0ns 0V 356240000.0ns 0V 356280000.0ns 0V 357080000.0ns 0V 357120000.0ns 0V 357840000.0ns 0V 357880000.0ns 0V 358360000.0ns 0V 358400000.0ns 0V 359120000.0ns 0V 359160000.0ns 0V 359960000.0ns 0V 360000000.0ns 0V 360080000.0ns 0V 360120000.0ns 0V 360920000.0ns 0V 360960000.0ns 0V 361680000.0ns 0V 361720000.0ns 0V 362200000.0ns 0V 362240000.0ns 0V 362960000.0ns 0V 363000000.0ns 0V 363800000.0ns 0V 363840000.0ns 0V 363920000.0ns 0V 363960000.0ns 0V 364760000.0ns 0V 364800000.0ns 0V 365520000.0ns 0V 365560000.0ns 0V 366040000.0ns 0V 366080000.0ns 0V 366800000.0ns 0V 366840000.0ns 0V 367640000.0ns 0V 367680000.0ns 0V 367760000.0ns 0V 367800000.0ns 0V 368600000.0ns 0V 368640000.0ns 0V 369360000.0ns 0V 369400000.0ns 0V 369880000.0ns 0V 369920000.0ns 0V 370640000.0ns 0V 370680000.0ns 0V 371480000.0ns 0V 371520000.0ns 0V 371600000.0ns 0V 371640000.0ns 0V 372440000.0ns 0V 372480000.0ns 0V 373200000.0ns 0V 373240000.0ns 0V 373720000.0ns 0V 373760000.0ns 0V 374480000.0ns 0V 374520000.0ns 0V 375320000.0ns 0V 375360000.0ns 0V 375440000.0ns 0V 375480000.0ns 0V 376280000.0ns 0V 376320000.0ns 0V 377040000.0ns 0V 377080000.0ns 0V 377560000.0ns 0V 377600000.0ns 0V 378320000.0ns 0V 378360000.0ns 0V 379160000.0ns 0V 379200000.0ns 0V 379280000.0ns 0V 379320000.0ns 0V 380120000.0ns 0V 380160000.0ns 0V 380880000.0ns 0V 380920000.0ns 0V 381400000.0ns 0V 381440000.0ns 0V 382160000.0ns 0V 382200000.0ns 0V 383000000.0ns 0V 383040000.0ns 0V 383120000.0ns 0V 383160000.0ns 0V 383960000.0ns 0V 384000000.0ns 0V 384720000.0ns 0V 384760000.0ns 0V 385240000.0ns 0V 385280000.0ns 0V 386000000.0ns 0V 386040000.0ns 0V 386840000.0ns 0V 386880000.0ns 0V 386960000.0ns 0V 387000000.0ns 0V 387800000.0ns 0V 387840000.0ns 0V 388560000.0ns 0V 388600000.0ns 0V 389080000.0ns 0V 389120000.0ns 0V 389840000.0ns 0V 389880000.0ns 0V 390680000.0ns 0V 390720000.0ns 0V 390800000.0ns 0V 390840000.0ns 0V)
VVWWL_J2 WWL_J2 0 PWL(0ns 0V 1800000.0ns 0V 1840000.0ns 1.95V 2240000.0ns 1.95V 2280000.0ns 0V 3960000.0ns 0V 7640000.0ns 0V 7680000.0ns 0V 8400000.0ns 0V 8440000.0ns 0V 8920000.0ns 0V 8960000.0ns 0V 9680000.0ns 0V 9720000.0ns 0V 10520000.0ns 0V 10560000.0ns 0V 10640000.0ns 0V 10680000.0ns 0V 11480000.0ns 0V 11520000.0ns 0V 12240000.0ns 0V 12280000.0ns 0V 12760000.0ns 0V 12800000.0ns 0V 13520000.0ns 0V 13560000.0ns 0V 14360000.0ns 0V 14400000.0ns 0V 14480000.0ns 0V 14520000.0ns 0V 15320000.0ns 0V 15360000.0ns 0V 16080000.0ns 0V 16120000.0ns 0V 16600000.0ns 0V 16640000.0ns 0V 17360000.0ns 0V 17400000.0ns 0V 18200000.0ns 0V 18240000.0ns 0V 18320000.0ns 0V 18360000.0ns 0V 19160000.0ns 0V 19200000.0ns 0V 19920000.0ns 0V 19960000.0ns 0V 20440000.0ns 0V 20480000.0ns 0V 21200000.0ns 0V 21240000.0ns 0V 22040000.0ns 0V 22080000.0ns 0V 22160000.0ns 0V 22200000.0ns 0V 23000000.0ns 0V 23040000.0ns 0V 23760000.0ns 0V 23800000.0ns 0V 24280000.0ns 0V 24320000.0ns 0V 25040000.0ns 0V 25080000.0ns 0V 25880000.0ns 0V 25920000.0ns 0V 26000000.0ns 0V 26040000.0ns 0V 26840000.0ns 0V 26880000.0ns 0V 27600000.0ns 0V 27640000.0ns 0V 28120000.0ns 0V 28160000.0ns 0V 28880000.0ns 0V 28920000.0ns 0V 29720000.0ns 0V 29760000.0ns 0V 29840000.0ns 0V 29880000.0ns 0V 30680000.0ns 0V 30720000.0ns 0V 31440000.0ns 0V 31480000.0ns 0V 31960000.0ns 0V 32000000.0ns 0V 32720000.0ns 0V 32760000.0ns 0V 33560000.0ns 0V 33600000.0ns 0V 33680000.0ns 0V 33720000.0ns 0V 34520000.0ns 0V 34560000.0ns 0V 35280000.0ns 0V 35320000.0ns 0V 35800000.0ns 0V 35840000.0ns 0V 36560000.0ns 0V 36600000.0ns 0V 37400000.0ns 0V 37440000.0ns 0V 37520000.0ns 0V 37560000.0ns 0V 38360000.0ns 0V 38400000.0ns 0V 39120000.0ns 0V 39160000.0ns 0V 39640000.0ns 0V 39680000.0ns 0V 40400000.0ns 0V 40440000.0ns 0V 41240000.0ns 0V 41280000.0ns 0V 41360000.0ns 0V 41400000.0ns 0V 42200000.0ns 0V 42240000.0ns 0V 42960000.0ns 0V 43000000.0ns 0V 43480000.0ns 0V 43520000.0ns 0V 44240000.0ns 0V 44280000.0ns 0V 45080000.0ns 0V 45120000.0ns 0V 45200000.0ns 0V 45240000.0ns 0V 46040000.0ns 0V 46080000.0ns 0V 46800000.0ns 0V 46840000.0ns 0V 47320000.0ns 0V 47360000.0ns 0V 48080000.0ns 0V 48120000.0ns 0V 48920000.0ns 0V 48960000.0ns 0V 49040000.0ns 0V 49080000.0ns 0V 49880000.0ns 0V 49920000.0ns 0V 50640000.0ns 0V 50680000.0ns 0V 51160000.0ns 0V 51200000.0ns 0V 51920000.0ns 0V 51960000.0ns 0V 52760000.0ns 0V 52800000.0ns 0V 52880000.0ns 0V 52920000.0ns 0V 53720000.0ns 0V 53760000.0ns 0V 54480000.0ns 0V 54520000.0ns 0V 55000000.0ns 0V 55040000.0ns 0V 55760000.0ns 0V 55800000.0ns 0V 56600000.0ns 0V 56640000.0ns 0V 56720000.0ns 0V 56760000.0ns 0V 57560000.0ns 0V 57600000.0ns 0V 58320000.0ns 0V 58360000.0ns 0V 58840000.0ns 0V 58880000.0ns 0V 59600000.0ns 0V 59640000.0ns 0V 60440000.0ns 0V 60480000.0ns 0V 60560000.0ns 0V 60600000.0ns 0V 61400000.0ns 0V 61440000.0ns 0V 62160000.0ns 0V 62200000.0ns 0V 62680000.0ns 0V 62720000.0ns 0V 63440000.0ns 0V 63480000.0ns 0V 64280000.0ns 0V 64320000.0ns 0V 64400000.0ns 0V 64440000.0ns 0V 65240000.0ns 0V 65280000.0ns 0V 66000000.0ns 0V 66040000.0ns 0V 66520000.0ns 0V 66560000.0ns 0V 67280000.0ns 0V 67320000.0ns 0V 68120000.0ns 0V 68160000.0ns 0V 68240000.0ns 0V 68280000.0ns 0V 69080000.0ns 0V 69120000.0ns 0V 69840000.0ns 0V 69880000.0ns 0V 70360000.0ns 0V 70400000.0ns 0V 71120000.0ns 0V 71160000.0ns 0V 71960000.0ns 0V 72000000.0ns 0V 72080000.0ns 0V 72120000.0ns 0V 72920000.0ns 0V 72960000.0ns 0V 73680000.0ns 0V 73720000.0ns 0V 74200000.0ns 0V 74240000.0ns 0V 74960000.0ns 0V 75000000.0ns 0V 75800000.0ns 0V 75840000.0ns 0V 75920000.0ns 0V 75960000.0ns 0V 76760000.0ns 0V 76800000.0ns 0V 77520000.0ns 0V 77560000.0ns 0V 78040000.0ns 0V 78080000.0ns 0V 78800000.0ns 0V 78840000.0ns 0V 79640000.0ns 0V 79680000.0ns 0V 79760000.0ns 0V 79800000.0ns 0V 80600000.0ns 0V 80640000.0ns 0V 81360000.0ns 0V 81400000.0ns 0V 81880000.0ns 0V 81920000.0ns 0V 82640000.0ns 0V 82680000.0ns 0V 83480000.0ns 0V 83520000.0ns 0V 83600000.0ns 0V 83640000.0ns 0V 84440000.0ns 0V 84480000.0ns 0V 85200000.0ns 0V 85240000.0ns 0V 85720000.0ns 0V 85760000.0ns 0V 86480000.0ns 0V 86520000.0ns 0V 87320000.0ns 0V 87360000.0ns 0V 87440000.0ns 0V 87480000.0ns 0V 88280000.0ns 0V 88320000.0ns 0V 89040000.0ns 0V 89080000.0ns 0V 89560000.0ns 0V 89600000.0ns 0V 90320000.0ns 0V 90360000.0ns 0V 91160000.0ns 0V 91200000.0ns 0V 91280000.0ns 0V 91320000.0ns 0V 92120000.0ns 0V 92160000.0ns 0V 92880000.0ns 0V 92920000.0ns 0V 93400000.0ns 0V 93440000.0ns 0V 94160000.0ns 0V 94200000.0ns 0V 95000000.0ns 0V 95040000.0ns 0V 95120000.0ns 0V 95160000.0ns 0V 95960000.0ns 0V 96000000.0ns 0V 96720000.0ns 0V 96760000.0ns 0V 97240000.0ns 0V 97280000.0ns 0V 98000000.0ns 0V 98040000.0ns 0V 98840000.0ns 0V 98880000.0ns 0V 98960000.0ns 0V 99000000.0ns 0V 99800000.0ns 0V 99840000.0ns 0V 100560000.0ns 0V 100600000.0ns 0V 101080000.0ns 0V 101120000.0ns 0V 101840000.0ns 0V 101880000.0ns 0V 102680000.0ns 0V 102720000.0ns 0V 102800000.0ns 0V 102840000.0ns 0V 103640000.0ns 0V 103680000.0ns 0V 104400000.0ns 0V 104440000.0ns 0V 104920000.0ns 0V 104960000.0ns 0V 105680000.0ns 0V 105720000.0ns 0V 106520000.0ns 0V 106560000.0ns 0V 106640000.0ns 0V 106680000.0ns 0V 107480000.0ns 0V 107520000.0ns 0V 108240000.0ns 0V 108280000.0ns 0V 108760000.0ns 0V 108800000.0ns 0V 109520000.0ns 0V 109560000.0ns 0V 110360000.0ns 0V 110400000.0ns 0V 110480000.0ns 0V 110520000.0ns 0V 111320000.0ns 0V 111360000.0ns 0V 112080000.0ns 0V 112120000.0ns 0V 112600000.0ns 0V 112640000.0ns 0V 113360000.0ns 0V 113400000.0ns 0V 114200000.0ns 0V 114240000.0ns 0V 114320000.0ns 0V 114360000.0ns 0V 115160000.0ns 0V 115200000.0ns 0V 115920000.0ns 0V 115960000.0ns 0V 116440000.0ns 0V 116480000.0ns 0V 117200000.0ns 0V 117240000.0ns 0V 118040000.0ns 0V 118080000.0ns 0V 118160000.0ns 0V 118200000.0ns 0V 119000000.0ns 0V 119040000.0ns 0V 119760000.0ns 0V 119800000.0ns 0V 120280000.0ns 0V 120320000.0ns 0V 121040000.0ns 0V 121080000.0ns 0V 121880000.0ns 0V 121920000.0ns 0V 122000000.0ns 0V 122040000.0ns 0V 122840000.0ns 0V 122880000.0ns 0V 123600000.0ns 0V 123640000.0ns 0V 124120000.0ns 0V 124160000.0ns 0V 124880000.0ns 0V 124920000.0ns 0V 125720000.0ns 0V 125760000.0ns 0V 125840000.0ns 0V 125880000.0ns 0V 126680000.0ns 0V 126720000.0ns 0V 127440000.0ns 0V 127480000.0ns 0V 127960000.0ns 0V 128000000.0ns 0V 128720000.0ns 0V 128760000.0ns 0V 129560000.0ns 0V 129600000.0ns 0V 129680000.0ns 0V 129720000.0ns 0V 130520000.0ns 0V 130560000.0ns 0V 131280000.0ns 0V 131320000.0ns 0V 131800000.0ns 0V 131840000.0ns 0V 132560000.0ns 0V 132600000.0ns 0V 133400000.0ns 0V 133440000.0ns 0V 133520000.0ns 0V 133560000.0ns 0V 134360000.0ns 0V 134400000.0ns 0V 135120000.0ns 0V 135160000.0ns 0V 135640000.0ns 0V 135680000.0ns 0V 136400000.0ns 0V 136440000.0ns 0V 137240000.0ns 0V 137280000.0ns 0V 137360000.0ns 0V 137400000.0ns 0V 138200000.0ns 0V 138240000.0ns 0V 138960000.0ns 0V 139000000.0ns 0V 139480000.0ns 0V 139520000.0ns 0V 140240000.0ns 0V 140280000.0ns 0V 141080000.0ns 0V 141120000.0ns 0V 141200000.0ns 0V 141240000.0ns 0V 142040000.0ns 0V 142080000.0ns 0V 142800000.0ns 0V 142840000.0ns 0V 143320000.0ns 0V 143360000.0ns 0V 144080000.0ns 0V 144120000.0ns 0V 144920000.0ns 0V 144960000.0ns 0V 145040000.0ns 0V 145080000.0ns 0V 145880000.0ns 0V 145920000.0ns 0V 146640000.0ns 0V 146680000.0ns 0V 147160000.0ns 0V 147200000.0ns 0V 147920000.0ns 0V 147960000.0ns 0V 148760000.0ns 0V 148800000.0ns 0V 148880000.0ns 0V 148920000.0ns 0V 149720000.0ns 0V 149760000.0ns 0V 150480000.0ns 0V 150520000.0ns 0V 151000000.0ns 0V 151040000.0ns 0V 151760000.0ns 0V 151800000.0ns 0V 152600000.0ns 0V 152640000.0ns 0V 152720000.0ns 0V 152760000.0ns 0V 153560000.0ns 0V 153600000.0ns 0V 154320000.0ns 0V 154360000.0ns 0V 154840000.0ns 0V 154880000.0ns 0V 155600000.0ns 0V 155640000.0ns 0V 156440000.0ns 0V 156480000.0ns 0V 156560000.0ns 0V 156600000.0ns 0V 157400000.0ns 0V 157440000.0ns 0V 158160000.0ns 0V 158200000.0ns 0V 158680000.0ns 0V 158720000.0ns 0V 159440000.0ns 0V 159480000.0ns 0V 160280000.0ns 0V 160320000.0ns 0V 160400000.0ns 0V 160440000.0ns 0V 161240000.0ns 0V 161280000.0ns 0V 162000000.0ns 0V 162040000.0ns 0V 162520000.0ns 0V 162560000.0ns 0V 163280000.0ns 0V 163320000.0ns 0V 164120000.0ns 0V 164160000.0ns 0V 164240000.0ns 0V 164280000.0ns 0V 165080000.0ns 0V 165120000.0ns 0V 165840000.0ns 0V 165880000.0ns 0V 166360000.0ns 0V 166400000.0ns 0V 167120000.0ns 0V 167160000.0ns 0V 167960000.0ns 0V 168000000.0ns 0V 168080000.0ns 0V 168120000.0ns 0V 168920000.0ns 0V 168960000.0ns 0V 169680000.0ns 0V 169720000.0ns 0V 170200000.0ns 0V 170240000.0ns 0V 170960000.0ns 0V 171000000.0ns 0V 171800000.0ns 0V 171840000.0ns 0V 171920000.0ns 0V 171960000.0ns 0V 172760000.0ns 0V 172800000.0ns 0V 173520000.0ns 0V 173560000.0ns 0V 174040000.0ns 0V 174080000.0ns 0V 174800000.0ns 0V 174840000.0ns 0V 175640000.0ns 0V 175680000.0ns 0V 175760000.0ns 0V 175800000.0ns 0V 176600000.0ns 0V 176640000.0ns 0V 177360000.0ns 0V 177400000.0ns 0V 177880000.0ns 0V 177920000.0ns 0V 178640000.0ns 0V 178680000.0ns 0V 179480000.0ns 0V 179520000.0ns 0V 179600000.0ns 0V 179640000.0ns 0V 180440000.0ns 0V 180480000.0ns 0V 181200000.0ns 0V 181240000.0ns 0V 181720000.0ns 0V 181760000.0ns 0V 182480000.0ns 0V 182520000.0ns 0V 183320000.0ns 0V 183360000.0ns 0V 183440000.0ns 0V 183480000.0ns 0V 184280000.0ns 0V 184320000.0ns 0V 185040000.0ns 0V 185080000.0ns 0V 185560000.0ns 0V 185600000.0ns 0V 186320000.0ns 0V 186360000.0ns 0V 187160000.0ns 0V 187200000.0ns 0V 187280000.0ns 0V 187320000.0ns 0V 188120000.0ns 0V 188160000.0ns 0V 188880000.0ns 0V 188920000.0ns 0V 189400000.0ns 0V 189440000.0ns 0V 190160000.0ns 0V 190200000.0ns 0V 191000000.0ns 0V 191040000.0ns 0V 191120000.0ns 0V 191160000.0ns 0V 191960000.0ns 0V 192000000.0ns 0V 192720000.0ns 0V 192760000.0ns 0V 193240000.0ns 0V 193280000.0ns 0V 194000000.0ns 0V 194040000.0ns 0V 194840000.0ns 0V 194880000.0ns 0V 194960000.0ns 0V 195000000.0ns 0V 195800000.0ns 0V 195840000.0ns 0V 196560000.0ns 0V 196600000.0ns 0V 197080000.0ns 0V 197120000.0ns 0V 197840000.0ns 0V 197880000.0ns 0V 198680000.0ns 0V 198720000.0ns 0V 198800000.0ns 0V 198840000.0ns 0V 199640000.0ns 0V 199680000.0ns 0V 200400000.0ns 0V 200440000.0ns 0V 200920000.0ns 0V 200960000.0ns 0V 201680000.0ns 0V 201720000.0ns 0V 202520000.0ns 0V 202560000.0ns 0V 202640000.0ns 0V 202680000.0ns 0V 203480000.0ns 0V 203520000.0ns 0V 204240000.0ns 0V 204280000.0ns 0V 204760000.0ns 0V 204800000.0ns 0V 205520000.0ns 0V 205560000.0ns 0V 206360000.0ns 0V 206400000.0ns 0V 206480000.0ns 0V 206520000.0ns 0V 207320000.0ns 0V 207360000.0ns 0V 208080000.0ns 0V 208120000.0ns 0V 208600000.0ns 0V 208640000.0ns 0V 209360000.0ns 0V 209400000.0ns 0V 210200000.0ns 0V 210240000.0ns 0V 210320000.0ns 0V 210360000.0ns 0V 211160000.0ns 0V 211200000.0ns 0V 211920000.0ns 0V 211960000.0ns 0V 212440000.0ns 0V 212480000.0ns 0V 213200000.0ns 0V 213240000.0ns 0V 214040000.0ns 0V 214080000.0ns 0V 214160000.0ns 0V 214200000.0ns 0V 215000000.0ns 0V 215040000.0ns 0V 215760000.0ns 0V 215800000.0ns 0V 216280000.0ns 0V 216320000.0ns 0V 217040000.0ns 0V 217080000.0ns 0V 217880000.0ns 0V 217920000.0ns 0V 218000000.0ns 0V 218040000.0ns 0V 218840000.0ns 0V 218880000.0ns 0V 219600000.0ns 0V 219640000.0ns 0V 220120000.0ns 0V 220160000.0ns 0V 220880000.0ns 0V 220920000.0ns 0V 221720000.0ns 0V 221760000.0ns 0V 221840000.0ns 0V 221880000.0ns 0V 222680000.0ns 0V 222720000.0ns 0V 223440000.0ns 0V 223480000.0ns 0V 223960000.0ns 0V 224000000.0ns 0V 224720000.0ns 0V 224760000.0ns 0V 225560000.0ns 0V 225600000.0ns 0V 225680000.0ns 0V 225720000.0ns 0V 226520000.0ns 0V 226560000.0ns 0V 227280000.0ns 0V 227320000.0ns 0V 227800000.0ns 0V 227840000.0ns 0V 228560000.0ns 0V 228600000.0ns 0V 229400000.0ns 0V 229440000.0ns 0V 229520000.0ns 0V 229560000.0ns 0V 230360000.0ns 0V 230400000.0ns 0V 231120000.0ns 0V 231160000.0ns 0V 231640000.0ns 0V 231680000.0ns 0V 232400000.0ns 0V 232440000.0ns 0V 233240000.0ns 0V 233280000.0ns 0V 233360000.0ns 0V 233400000.0ns 0V 234200000.0ns 0V 234240000.0ns 0V 234960000.0ns 0V 235000000.0ns 0V 235480000.0ns 0V 235520000.0ns 0V 236240000.0ns 0V 236280000.0ns 0V 237080000.0ns 0V 237120000.0ns 0V 237200000.0ns 0V 237240000.0ns 0V 238040000.0ns 0V 238080000.0ns 0V 238800000.0ns 0V 238840000.0ns 0V 239320000.0ns 0V 239360000.0ns 0V 240080000.0ns 0V 240120000.0ns 0V 240920000.0ns 0V 240960000.0ns 0V 241040000.0ns 0V 241080000.0ns 0V 241880000.0ns 0V 241920000.0ns 0V 242640000.0ns 0V 242680000.0ns 0V 243160000.0ns 0V 243200000.0ns 0V 243920000.0ns 0V 243960000.0ns 0V 244760000.0ns 0V 244800000.0ns 0V 244880000.0ns 0V 244920000.0ns 0V 245720000.0ns 0V 245760000.0ns 0V 246480000.0ns 0V 246520000.0ns 0V 247000000.0ns 0V 247040000.0ns 0V 247760000.0ns 0V 247800000.0ns 0V 248600000.0ns 0V 248640000.0ns 0V 248720000.0ns 0V 248760000.0ns 0V 249560000.0ns 0V 249600000.0ns 0V 250320000.0ns 0V 250360000.0ns 0V 250840000.0ns 0V 250880000.0ns 0V 251600000.0ns 0V 251640000.0ns 0V 252440000.0ns 0V 252480000.0ns 0V 252560000.0ns 0V 252600000.0ns 0V 253400000.0ns 0V 253440000.0ns 0V 254160000.0ns 0V 254200000.0ns 0V 254680000.0ns 0V 254720000.0ns 0V 255440000.0ns 0V 255480000.0ns 0V 256280000.0ns 0V 256320000.0ns 0V 256400000.0ns 0V 256440000.0ns 0V 257240000.0ns 0V 257280000.0ns 0V 258000000.0ns 0V 258040000.0ns 0V 258520000.0ns 0V 258560000.0ns 0V 259280000.0ns 0V 259320000.0ns 0V 260120000.0ns 0V 260160000.0ns 0V 260240000.0ns 0V 260280000.0ns 0V 261080000.0ns 0V 261120000.0ns 0V 261840000.0ns 0V 261880000.0ns 0V 262360000.0ns 0V 262400000.0ns 0V 263120000.0ns 0V 263160000.0ns 0V 263960000.0ns 0V 264000000.0ns 0V 264080000.0ns 0V 264120000.0ns 0V 264920000.0ns 0V 264960000.0ns 0V 265680000.0ns 0V 265720000.0ns 0V 266200000.0ns 0V 266240000.0ns 0V 266960000.0ns 0V 267000000.0ns 0V 267800000.0ns 0V 267840000.0ns 0V 267920000.0ns 0V 267960000.0ns 0V 268760000.0ns 0V 268800000.0ns 0V 269520000.0ns 0V 269560000.0ns 0V 270040000.0ns 0V 270080000.0ns 0V 270800000.0ns 0V 270840000.0ns 0V 271640000.0ns 0V 271680000.0ns 0V 271760000.0ns 0V 271800000.0ns 0V 272600000.0ns 0V 272640000.0ns 0V 273360000.0ns 0V 273400000.0ns 0V 273880000.0ns 0V 273920000.0ns 0V 274640000.0ns 0V 274680000.0ns 0V 275480000.0ns 0V 275520000.0ns 0V 275600000.0ns 0V 275640000.0ns 0V 276440000.0ns 0V 276480000.0ns 0V 277200000.0ns 0V 277240000.0ns 0V 277720000.0ns 0V 277760000.0ns 0V 278480000.0ns 0V 278520000.0ns 0V 279320000.0ns 0V 279360000.0ns 0V 279440000.0ns 0V 279480000.0ns 0V 280280000.0ns 0V 280320000.0ns 0V 281040000.0ns 0V 281080000.0ns 0V 281560000.0ns 0V 281600000.0ns 0V 282320000.0ns 0V 282360000.0ns 0V 283160000.0ns 0V 283200000.0ns 0V 283280000.0ns 0V 283320000.0ns 0V 284120000.0ns 0V 284160000.0ns 0V 284880000.0ns 0V 284920000.0ns 0V 285400000.0ns 0V 285440000.0ns 0V 286160000.0ns 0V 286200000.0ns 0V 287000000.0ns 0V 287040000.0ns 0V 287120000.0ns 0V 287160000.0ns 0V 287960000.0ns 0V 288000000.0ns 0V 288720000.0ns 0V 288760000.0ns 0V 289240000.0ns 0V 289280000.0ns 0V 290000000.0ns 0V 290040000.0ns 0V 290840000.0ns 0V 290880000.0ns 0V 290960000.0ns 0V 291000000.0ns 0V 291800000.0ns 0V 291840000.0ns 0V 292560000.0ns 0V 292600000.0ns 0V 293080000.0ns 0V 293120000.0ns 0V 293840000.0ns 0V 293880000.0ns 0V 294680000.0ns 0V 294720000.0ns 0V 294800000.0ns 0V 294840000.0ns 0V 295640000.0ns 0V 295680000.0ns 0V 296400000.0ns 0V 296440000.0ns 0V 296920000.0ns 0V 296960000.0ns 0V 297680000.0ns 0V 297720000.0ns 0V 298520000.0ns 0V 298560000.0ns 0V 298640000.0ns 0V 298680000.0ns 0V 299480000.0ns 0V 299520000.0ns 0V 300240000.0ns 0V 300280000.0ns 0V 300760000.0ns 0V 300800000.0ns 0V 301520000.0ns 0V 301560000.0ns 0V 302360000.0ns 0V 302400000.0ns 0V 302480000.0ns 0V 302520000.0ns 0V 303320000.0ns 0V 303360000.0ns 0V 304080000.0ns 0V 304120000.0ns 0V 304600000.0ns 0V 304640000.0ns 0V 305360000.0ns 0V 305400000.0ns 0V 306200000.0ns 0V 306240000.0ns 0V 306320000.0ns 0V 306360000.0ns 0V 307160000.0ns 0V 307200000.0ns 0V 307920000.0ns 0V 307960000.0ns 0V 308440000.0ns 0V 308480000.0ns 0V 309200000.0ns 0V 309240000.0ns 0V 310040000.0ns 0V 310080000.0ns 0V 310160000.0ns 0V 310200000.0ns 0V 311000000.0ns 0V 311040000.0ns 0V 311760000.0ns 0V 311800000.0ns 0V 312280000.0ns 0V 312320000.0ns 0V 313040000.0ns 0V 313080000.0ns 0V 313880000.0ns 0V 313920000.0ns 0V 314000000.0ns 0V 314040000.0ns 0V 314840000.0ns 0V 314880000.0ns 0V 315600000.0ns 0V 315640000.0ns 0V 316120000.0ns 0V 316160000.0ns 0V 316880000.0ns 0V 316920000.0ns 0V 317720000.0ns 0V 317760000.0ns 0V 317840000.0ns 0V 317880000.0ns 0V 318680000.0ns 0V 318720000.0ns 0V 319440000.0ns 0V 319480000.0ns 0V 319960000.0ns 0V 320000000.0ns 0V 320720000.0ns 0V 320760000.0ns 0V 321560000.0ns 0V 321600000.0ns 0V 321680000.0ns 0V 321720000.0ns 0V 322520000.0ns 0V 322560000.0ns 0V 323280000.0ns 0V 323320000.0ns 0V 323800000.0ns 0V 323840000.0ns 0V 324560000.0ns 0V 324600000.0ns 0V 325400000.0ns 0V 325440000.0ns 0V 325520000.0ns 0V 325560000.0ns 0V 326360000.0ns 0V 326400000.0ns 0V 327120000.0ns 0V 327160000.0ns 0V 327640000.0ns 0V 327680000.0ns 0V 328400000.0ns 0V 328440000.0ns 0V 329240000.0ns 0V 329280000.0ns 0V 329360000.0ns 0V 329400000.0ns 0V 330200000.0ns 0V 330240000.0ns 0V 330960000.0ns 0V 331000000.0ns 0V 331480000.0ns 0V 331520000.0ns 0V 332240000.0ns 0V 332280000.0ns 0V 333080000.0ns 0V 333120000.0ns 0V 333200000.0ns 0V 333240000.0ns 0V 334040000.0ns 0V 334080000.0ns 0V 334800000.0ns 0V 334840000.0ns 0V 335320000.0ns 0V 335360000.0ns 0V 336080000.0ns 0V 336120000.0ns 0V 336920000.0ns 0V 336960000.0ns 0V 337040000.0ns 0V 337080000.0ns 0V 337880000.0ns 0V 337920000.0ns 0V 338640000.0ns 0V 338680000.0ns 0V 339160000.0ns 0V 339200000.0ns 0V 339920000.0ns 0V 339960000.0ns 0V 340760000.0ns 0V 340800000.0ns 0V 340880000.0ns 0V 340920000.0ns 0V 341720000.0ns 0V 341760000.0ns 0V 342480000.0ns 0V 342520000.0ns 0V 343000000.0ns 0V 343040000.0ns 0V 343760000.0ns 0V 343800000.0ns 0V 344600000.0ns 0V 344640000.0ns 0V 344720000.0ns 0V 344760000.0ns 0V 345560000.0ns 0V 345600000.0ns 0V 346320000.0ns 0V 346360000.0ns 0V 346840000.0ns 0V 346880000.0ns 0V 347600000.0ns 0V 347640000.0ns 0V 348440000.0ns 0V 348480000.0ns 0V 348560000.0ns 0V 348600000.0ns 0V 349400000.0ns 0V 349440000.0ns 0V 350160000.0ns 0V 350200000.0ns 0V 350680000.0ns 0V 350720000.0ns 0V 351440000.0ns 0V 351480000.0ns 0V 352280000.0ns 0V 352320000.0ns 0V 352400000.0ns 0V 352440000.0ns 0V 353240000.0ns 0V 353280000.0ns 0V 354000000.0ns 0V 354040000.0ns 0V 354520000.0ns 0V 354560000.0ns 0V 355280000.0ns 0V 355320000.0ns 0V 356120000.0ns 0V 356160000.0ns 0V 356240000.0ns 0V 356280000.0ns 0V 357080000.0ns 0V 357120000.0ns 0V 357840000.0ns 0V 357880000.0ns 0V 358360000.0ns 0V 358400000.0ns 0V 359120000.0ns 0V 359160000.0ns 0V 359960000.0ns 0V 360000000.0ns 0V 360080000.0ns 0V 360120000.0ns 0V 360920000.0ns 0V 360960000.0ns 0V 361680000.0ns 0V 361720000.0ns 0V 362200000.0ns 0V 362240000.0ns 0V 362960000.0ns 0V 363000000.0ns 0V 363800000.0ns 0V 363840000.0ns 0V 363920000.0ns 0V 363960000.0ns 0V 364760000.0ns 0V 364800000.0ns 0V 365520000.0ns 0V 365560000.0ns 0V 366040000.0ns 0V 366080000.0ns 0V 366800000.0ns 0V 366840000.0ns 0V 367640000.0ns 0V 367680000.0ns 0V 367760000.0ns 0V 367800000.0ns 0V 368600000.0ns 0V 368640000.0ns 0V 369360000.0ns 0V 369400000.0ns 0V 369880000.0ns 0V 369920000.0ns 0V 370640000.0ns 0V 370680000.0ns 0V 371480000.0ns 0V 371520000.0ns 0V 371600000.0ns 0V 371640000.0ns 0V 372440000.0ns 0V 372480000.0ns 0V 373200000.0ns 0V 373240000.0ns 0V 373720000.0ns 0V 373760000.0ns 0V 374480000.0ns 0V 374520000.0ns 0V 375320000.0ns 0V 375360000.0ns 0V 375440000.0ns 0V 375480000.0ns 0V 376280000.0ns 0V 376320000.0ns 0V 377040000.0ns 0V 377080000.0ns 0V 377560000.0ns 0V 377600000.0ns 0V 378320000.0ns 0V 378360000.0ns 0V 379160000.0ns 0V 379200000.0ns 0V 379280000.0ns 0V 379320000.0ns 0V 380120000.0ns 0V 380160000.0ns 0V 380880000.0ns 0V 380920000.0ns 0V 381400000.0ns 0V 381440000.0ns 0V 382160000.0ns 0V 382200000.0ns 0V 383000000.0ns 0V 383040000.0ns 0V 383120000.0ns 0V 383160000.0ns 0V 383960000.0ns 0V 384000000.0ns 0V 384720000.0ns 0V 384760000.0ns 0V 385240000.0ns 0V 385280000.0ns 0V 386000000.0ns 0V 386040000.0ns 0V 386840000.0ns 0V 386880000.0ns 0V 386960000.0ns 0V 387000000.0ns 0V 387800000.0ns 0V 387840000.0ns 0V 388560000.0ns 0V 388600000.0ns 0V 389080000.0ns 0V 389120000.0ns 0V 389840000.0ns 0V 389880000.0ns 0V 390680000.0ns 0V 390720000.0ns 0V 390800000.0ns 0V 390840000.0ns 0V)
.model switch VSWITCH (ROFF=100000000000.0kOhm RON=0.0001Ohm VOFF=0.4V VON=0.5V)
.model NMOSS NMOS (A0=1.5 A1=0.0 A2=0.42385546 AGS=1.25 ALPHA0=3e-08 ALPHA1=0.85 B0=0.0 B1=0.0 BETA0=13.85 CGBO=1e-13 CGDO=2.54e-10 CGSO=2.54e-10 DELTA=0.01 DR0UT=0.50332666 DVT0=0.0 DVT1=0.53 DVT2=-0.032 ETA0=0.00069413878 K1=0.90707349 K2=-0.12949 K3=2.0 KETA=0.0 L=0.15 LEVEL=54 LINT=1.1932e-08 NDEP=1.7e+17 NFACTOR=2.015 NSUB=1e+20 PCLM=0.14094 PDIBLC1=0.35697215 PDIBLC2=0.0084061121 PDIBLCB=-0.10329577 PRWB=0.0 PRWG=0.021507 PSCBE1=791419880.0 PSCBE2=1e-12 PVAG=0.0 RDSW=65.968 RSH=0.1 TOX=4.148e-09 U0=0.030197 VOFF=-0.20753 VSAT=176320 VTO=0.7 W=10 WINT=2.1859e-08 XJ=1.5e-07)
.model diode D ()
.model capacitor C ()
.ends mlp
Xmlp NUDGED FREE X_0 X_1 X_2 Y_0_NUDGED Y_1_NUDGED mlp
.options TEMP = 27
.options TNOM = 27
.tran 20000ns 474085920.0ns 0s
.end
